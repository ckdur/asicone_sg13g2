VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.34 BY 6.12 ;
END obssite

#--------EOF---------

MACRO AN2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1
MACRO AN2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 1.350 0.815 2.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 1.350 1.775 2.170 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 0.335 2.650 ;
        RECT 0.175 2.490 2.735 2.650 ;
        RECT 2.525 2.490 2.785 2.650 ;
  END
END AN2D1_1
MACRO AN2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1_2
MACRO AN2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 2.255 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1_3
#--------EOF---------

MACRO AN2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1
MACRO AN2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 1.350 0.815 2.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 1.350 1.775 2.170 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 0.335 2.650 ;
        RECT 0.175 2.490 2.735 2.650 ;
        RECT 2.525 2.490 2.785 2.650 ;
  END
END AN2D1_1
MACRO AN2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1_2
MACRO AN2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 2.255 1.110 ;
        RECT 2.095 0.950 2.255 3.610 ;
        RECT 2.045 3.450 2.305 3.610 ;
  END
END AN2D1_3
#--------EOF---------

MACRO AO21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 1.775 3.610 ;
        RECT 1.565 3.450 1.825 3.610 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 2.575 2.490 2.735 3.610 ;
        RECT 2.525 3.450 2.785 3.610 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 1.295 1.110 ;
        RECT 1.135 0.950 1.295 3.130 ;
        RECT 1.085 2.970 1.345 3.130 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 3.055 0.950 3.215 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.175 4.210 0.335 4.830 ;
        RECT 0.175 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END AO21D1
MACRO AO21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.525 4.670 2.785 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 2.575 0.950 3.215 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 3.055 4.210 3.215 4.830 ;
  END
END AO21D1_1
MACRO AO21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 1.135 0.290 4.655 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AO21D1_2
MACRO AO21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 0.175 5.010 2.255 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
  END
END AO21D1_3
#--------EOF---------

MACRO AO21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 1.775 3.610 ;
        RECT 1.565 3.450 1.825 3.610 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 2.575 2.490 2.735 3.610 ;
        RECT 2.525 3.450 2.785 3.610 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 1.295 1.110 ;
        RECT 1.135 0.950 1.295 3.130 ;
        RECT 1.085 2.970 1.345 3.130 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 3.055 0.950 3.215 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.175 4.210 0.335 4.830 ;
        RECT 0.175 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END AO21D1
MACRO AO21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.525 4.670 2.785 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 2.575 0.950 3.215 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 3.055 4.210 3.215 4.830 ;
  END
END AO21D1_1
MACRO AO21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 1.135 0.290 4.655 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AO21D1_2
MACRO AO21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 0.175 5.010 2.255 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
  END
END AO21D1_3
#--------EOF---------

MACRO AOI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 2.255 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
  END
END AOI21D1
MACRO AOI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 4.670 3.215 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 1.135 4.670 1.295 5.170 ;
  END
END AOI21D1_1
MACRO AOI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 2.010 0.385 2.170 ;
        RECT 0.175 2.010 0.335 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.655 0.950 2.255 1.110 ;
        RECT 0.655 0.950 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 0.655 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AOI21D1_2
MACRO AOI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.210 2.255 4.370 ;
        RECT 0.175 4.210 0.335 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AOI21D1_3
#--------EOF---------

MACRO AOI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 2.255 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
  END
END AOI21D1
MACRO AOI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 4.670 3.215 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 1.135 4.670 1.295 5.170 ;
  END
END AOI21D1_1
MACRO AOI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 2.010 0.385 2.170 ;
        RECT 0.175 2.010 0.335 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.655 0.950 2.255 1.110 ;
        RECT 0.655 0.950 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 0.655 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AOI21D1_2
MACRO AOI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.210 2.255 4.370 ;
        RECT 0.175 4.210 0.335 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 4.670 1.295 5.170 ;
        RECT 1.135 5.010 3.215 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
  END
END AOI21D1_3
#--------EOF---------

MACRO BUFFD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 1.775 3.610 ;
        RECT 1.615 3.450 1.775 5.170 ;
        RECT 1.615 5.010 2.255 5.170 ;
        RECT 0.655 0.950 2.255 1.110 ;
        RECT 0.655 0.950 0.815 2.170 ;
        RECT 0.605 2.010 0.865 2.170 ;
  END
END BUFFD1
MACRO BUFFD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 0.655 3.450 1.775 3.610 ;
        RECT 0.655 3.450 0.815 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.950 1.775 2.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
  END
END BUFFD1_1
#--------EOF---------

MACRO BUFFD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 1.775 3.610 ;
        RECT 1.615 3.450 1.775 5.170 ;
        RECT 1.615 5.010 2.255 5.170 ;
        RECT 0.655 0.950 2.255 1.110 ;
        RECT 0.655 0.950 0.815 2.170 ;
        RECT 0.605 2.010 0.865 2.170 ;
  END
END BUFFD1
MACRO BUFFD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 0.655 3.450 1.775 3.610 ;
        RECT 0.655 3.450 0.815 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.950 1.775 2.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
  END
END BUFFD1_1
#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFCNQD1 0 0 ; 
  SIZE 17.000 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cdn
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 7.375 2.010 8.015 2.170 ;
    END 
  END cdn
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 16.445 0.950 16.705 1.110 ;
        RECT 15.485 4.670 15.745 4.830 ;
        RECT 16.495 0.950 16.655 4.370 ;
        RECT 15.535 4.210 16.655 4.370 ;
        RECT 15.535 4.210 15.695 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 8.765 5.010 9.025 5.170 ;
        RECT 8.815 5.010 8.975 6.050 ;
        RECT 12.605 5.010 12.865 5.170 ;
        RECT 12.655 5.010 12.815 6.050 ;
        RECT 0.000 6.020 17.000 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.855 0.070 8.015 1.110 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.655 0.070 12.815 1.110 ;
        RECT 15.485 0.950 15.745 1.110 ;
        RECT 15.535 0.070 15.695 1.110 ;
        RECT 0.000 -0.100 17.000 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.290 1.775 1.110 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 10.415 3.130 ;
        RECT 10.205 2.970 10.465 3.130 ;
        RECT 0.175 5.010 0.335 5.830 ;
        RECT 0.175 5.670 1.775 5.830 ;
        RECT 1.565 5.670 1.825 5.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 5.170 ;
        RECT 2.045 4.210 2.305 4.370 ;
        RECT 2.095 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 3.535 3.450 5.615 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
        RECT 8.765 3.450 9.025 3.610 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 2.650 ;
        RECT 4.975 2.490 9.455 2.650 ;
        RECT 9.245 2.490 9.505 2.650 ;
        RECT 8.285 2.490 8.545 2.650 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 4.975 4.210 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
        RECT 4.925 2.490 5.185 2.650 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 7.805 5.010 8.065 5.170 ;
        RECT 5.935 5.010 8.015 5.170 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 8.815 0.950 8.975 1.510 ;
        RECT 6.415 1.350 8.975 1.510 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.365 4.210 6.625 4.370 ;
        RECT 6.415 4.210 9.935 4.370 ;
        RECT 9.775 4.210 9.935 4.830 ;
        RECT 9.725 0.950 9.985 1.110 ;
        RECT 10.685 4.670 10.945 4.830 ;
        RECT 9.775 0.290 9.935 1.110 ;
        RECT 9.775 0.290 12.335 0.450 ;
        RECT 12.125 0.290 12.385 0.450 ;
        RECT 14.045 2.010 14.305 2.170 ;
        RECT 14.095 2.010 14.255 4.370 ;
        RECT 10.735 4.210 14.255 4.370 ;
        RECT 10.735 4.210 10.895 4.830 ;
        RECT 14.045 3.450 14.305 3.610 ;
        RECT 10.685 0.950 10.945 1.110 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.735 0.950 11.855 1.110 ;
        RECT 14.525 0.950 14.785 1.110 ;
        RECT 13.565 4.670 13.825 4.830 ;
        RECT 12.125 1.350 12.385 1.510 ;
        RECT 12.175 1.350 14.735 1.510 ;
        RECT 14.575 0.950 14.735 1.510 ;
        RECT 14.575 1.350 14.735 4.830 ;
        RECT 13.615 4.670 14.735 4.830 ;
  END
END DFCNQD1
#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFCNQD1 0 0 ; 
  SIZE 17.000 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cdn
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 7.375 2.010 8.015 2.170 ;
    END 
  END cdn
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 16.445 0.950 16.705 1.110 ;
        RECT 15.485 4.670 15.745 4.830 ;
        RECT 16.495 0.950 16.655 4.370 ;
        RECT 15.535 4.210 16.655 4.370 ;
        RECT 15.535 4.210 15.695 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 8.765 5.010 9.025 5.170 ;
        RECT 8.815 5.010 8.975 6.050 ;
        RECT 12.605 5.010 12.865 5.170 ;
        RECT 12.655 5.010 12.815 6.050 ;
        RECT 0.000 6.020 17.000 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.855 0.070 8.015 1.110 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.655 0.070 12.815 1.110 ;
        RECT 15.485 0.950 15.745 1.110 ;
        RECT 15.535 0.070 15.695 1.110 ;
        RECT 0.000 -0.100 17.000 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.290 1.775 1.110 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 10.415 3.130 ;
        RECT 10.205 2.970 10.465 3.130 ;
        RECT 0.175 5.010 0.335 5.830 ;
        RECT 0.175 5.670 1.775 5.830 ;
        RECT 1.565 5.670 1.825 5.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 5.170 ;
        RECT 2.045 4.210 2.305 4.370 ;
        RECT 2.095 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 3.535 3.450 5.615 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
        RECT 8.765 3.450 9.025 3.610 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 2.650 ;
        RECT 4.975 2.490 9.455 2.650 ;
        RECT 9.245 2.490 9.505 2.650 ;
        RECT 8.285 2.490 8.545 2.650 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 4.975 4.210 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
        RECT 4.925 2.490 5.185 2.650 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 7.805 5.010 8.065 5.170 ;
        RECT 5.935 5.010 8.015 5.170 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 8.815 0.950 8.975 1.510 ;
        RECT 6.415 1.350 8.975 1.510 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.365 4.210 6.625 4.370 ;
        RECT 6.415 4.210 9.935 4.370 ;
        RECT 9.775 4.210 9.935 4.830 ;
        RECT 9.725 0.950 9.985 1.110 ;
        RECT 10.685 4.670 10.945 4.830 ;
        RECT 9.775 0.290 9.935 1.110 ;
        RECT 9.775 0.290 12.335 0.450 ;
        RECT 12.125 0.290 12.385 0.450 ;
        RECT 14.045 2.010 14.305 2.170 ;
        RECT 14.095 2.010 14.255 4.370 ;
        RECT 10.735 4.210 14.255 4.370 ;
        RECT 10.735 4.210 10.895 4.830 ;
        RECT 14.045 3.450 14.305 3.610 ;
        RECT 10.685 0.950 10.945 1.110 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.735 0.950 11.855 1.110 ;
        RECT 14.525 0.950 14.785 1.110 ;
        RECT 13.565 4.670 13.825 4.830 ;
        RECT 12.125 1.350 12.385 1.510 ;
        RECT 12.175 1.350 14.735 1.510 ;
        RECT 14.575 0.950 14.735 1.510 ;
        RECT 14.575 1.350 14.735 4.830 ;
        RECT 13.615 4.670 14.735 4.830 ;
  END
END DFCNQD1
#--------EOF---------

MACRO DFQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1 0 0 ; 
  SIZE 14.960 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.490 0.865 2.650 ;
        RECT 0.655 2.490 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 13.565 0.950 13.825 1.110 ;
        RECT 13.565 4.670 13.825 4.830 ;
        RECT 13.615 0.950 13.775 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.960 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.960 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.125 2.970 0.385 3.130 ;
        RECT 0.175 2.970 0.335 4.830 ;
        RECT 12.125 0.290 12.385 0.450 ;
        RECT 7.855 0.290 12.335 0.450 ;
        RECT 7.805 0.290 8.065 0.450 ;
        RECT 0.175 0.950 0.335 3.130 ;
        RECT 0.175 2.970 0.335 4.370 ;
        RECT 0.175 4.210 3.215 4.370 ;
        RECT 3.005 4.210 3.265 4.370 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 4.015 3.450 5.615 3.610 ;
        RECT 4.015 3.450 4.175 4.370 ;
        RECT 3.965 4.210 4.225 4.370 ;
        RECT 5.405 5.670 5.665 5.830 ;
        RECT 3.535 5.670 5.615 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 12.605 5.010 12.865 5.170 ;
        RECT 10.735 0.950 12.815 1.110 ;
        RECT 10.735 0.950 10.895 1.510 ;
        RECT 6.895 1.350 10.895 1.510 ;
        RECT 6.895 0.950 7.055 1.510 ;
        RECT 9.295 1.350 9.455 3.610 ;
        RECT 9.245 3.450 9.505 3.610 ;
        RECT 9.245 2.010 9.505 2.170 ;
        RECT 9.295 2.010 9.455 4.830 ;
        RECT 9.295 4.670 12.815 4.830 ;
        RECT 12.655 4.670 12.815 5.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.055 2.010 8.495 2.170 ;
        RECT 8.285 2.010 8.545 2.170 ;
        RECT 8.285 2.970 8.545 3.130 ;
        RECT 3.535 2.970 8.495 3.130 ;
        RECT 3.535 2.970 3.695 4.830 ;
        RECT 3.055 4.670 3.695 4.830 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 3.485 1.350 3.745 1.510 ;
        RECT 3.535 1.350 6.095 1.510 ;
        RECT 5.935 0.950 6.095 1.510 ;
        RECT 6.365 4.670 6.625 4.830 ;
        RECT 5.935 4.670 6.575 4.830 ;
        RECT 5.935 1.350 6.575 1.510 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 4.670 6.575 5.830 ;
        RECT 6.415 5.670 12.335 5.830 ;
        RECT 12.125 5.670 12.385 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 7.535 0.450 ;
        RECT 7.375 0.290 7.535 1.110 ;
        RECT 7.375 0.950 8.015 1.110 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 4.495 4.210 8.015 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
        RECT 9.725 0.950 9.985 1.110 ;
        RECT 11.165 1.350 11.425 1.510 ;
        RECT 11.215 1.350 13.295 1.510 ;
        RECT 13.085 1.350 13.345 1.510 ;
        RECT 10.205 0.950 10.465 1.110 ;
        RECT 9.775 0.950 10.415 1.110 ;
  END
END DFQD1
MACRO DFQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_1 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 0.175 0.290 1.775 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 9.245 2.010 9.505 2.170 ;
        RECT 9.295 2.010 9.455 3.610 ;
        RECT 9.245 3.450 9.505 3.610 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 0.335 5.830 ;
        RECT 0.175 5.670 3.695 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.775 3.450 9.935 4.370 ;
        RECT 8.815 4.210 9.935 4.370 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 3.055 2.490 7.535 2.650 ;
        RECT 7.325 2.490 7.585 2.650 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 3.055 2.010 7.535 2.170 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 3.485 4.210 3.745 4.370 ;
        RECT 3.535 4.210 3.695 4.830 ;
        RECT 3.535 4.670 6.095 4.830 ;
        RECT 8.285 0.290 8.545 0.450 ;
        RECT 5.935 0.290 8.495 0.450 ;
        RECT 5.935 0.290 6.095 1.110 ;
        RECT 5.935 4.670 6.095 5.830 ;
        RECT 5.935 5.670 9.455 5.830 ;
        RECT 9.245 5.670 9.505 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 4.495 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 7.855 1.350 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_1
MACRO DFQD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_2 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.950 1.775 2.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.295 3.450 9.935 3.610 ;
        RECT 9.295 3.450 9.455 4.830 ;
        RECT 8.815 4.670 9.455 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 4.975 0.290 7.535 0.450 ;
        RECT 7.325 0.290 7.585 0.450 ;
        RECT 7.325 4.210 7.585 4.370 ;
        RECT 4.975 4.210 7.535 4.370 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 5.405 1.350 5.665 1.510 ;
        RECT 2.095 1.350 5.615 1.510 ;
        RECT 2.095 0.950 2.255 1.510 ;
        RECT 8.285 2.010 8.545 2.170 ;
        RECT 2.575 2.010 8.495 2.170 ;
        RECT 2.575 2.010 2.735 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 5.455 1.350 5.615 2.170 ;
        RECT 8.335 2.010 8.495 5.830 ;
        RECT 8.335 5.670 9.455 5.830 ;
        RECT 9.245 5.670 9.505 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 3.535 5.670 8.495 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 6.365 3.450 6.625 3.610 ;
        RECT 6.415 3.450 8.015 3.610 ;
        RECT 7.855 3.450 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_2
MACRO DFQD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_3 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 2.970 1.345 3.130 ;
        RECT 1.135 2.970 1.295 3.610 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 9.245 0.290 9.505 0.450 ;
        RECT 4.015 0.290 9.455 0.450 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 2.575 0.950 4.175 1.110 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 1.775 2.170 ;
        RECT 1.615 2.010 1.775 4.830 ;
        RECT 1.615 4.670 2.255 4.830 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 0.655 2.490 2.255 2.650 ;
        RECT 0.605 2.490 0.865 2.650 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.295 3.450 9.935 3.610 ;
        RECT 9.295 3.450 9.455 4.830 ;
        RECT 8.815 4.670 9.455 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 4.975 2.010 7.535 2.170 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.175 0.290 3.695 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 8.495 5.170 ;
        RECT 8.335 3.450 8.495 5.170 ;
        RECT 8.285 3.450 8.545 3.610 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 3.535 5.010 3.695 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 7.855 1.350 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_3
#--------EOF---------

MACRO DFQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1 0 0 ; 
  SIZE 14.960 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.490 0.865 2.650 ;
        RECT 0.655 2.490 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 13.565 0.950 13.825 1.110 ;
        RECT 13.565 4.670 13.825 4.830 ;
        RECT 13.615 0.950 13.775 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.960 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.960 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.125 2.970 0.385 3.130 ;
        RECT 0.175 2.970 0.335 4.830 ;
        RECT 12.125 0.290 12.385 0.450 ;
        RECT 7.855 0.290 12.335 0.450 ;
        RECT 7.805 0.290 8.065 0.450 ;
        RECT 0.175 0.950 0.335 3.130 ;
        RECT 0.175 2.970 0.335 4.370 ;
        RECT 0.175 4.210 3.215 4.370 ;
        RECT 3.005 4.210 3.265 4.370 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 4.015 3.450 5.615 3.610 ;
        RECT 4.015 3.450 4.175 4.370 ;
        RECT 3.965 4.210 4.225 4.370 ;
        RECT 5.405 5.670 5.665 5.830 ;
        RECT 3.535 5.670 5.615 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 12.605 5.010 12.865 5.170 ;
        RECT 10.735 0.950 12.815 1.110 ;
        RECT 10.735 0.950 10.895 1.510 ;
        RECT 6.895 1.350 10.895 1.510 ;
        RECT 6.895 0.950 7.055 1.510 ;
        RECT 9.295 1.350 9.455 3.610 ;
        RECT 9.245 3.450 9.505 3.610 ;
        RECT 9.245 2.010 9.505 2.170 ;
        RECT 9.295 2.010 9.455 4.830 ;
        RECT 9.295 4.670 12.815 4.830 ;
        RECT 12.655 4.670 12.815 5.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.055 2.010 8.495 2.170 ;
        RECT 8.285 2.010 8.545 2.170 ;
        RECT 8.285 2.970 8.545 3.130 ;
        RECT 3.535 2.970 8.495 3.130 ;
        RECT 3.535 2.970 3.695 4.830 ;
        RECT 3.055 4.670 3.695 4.830 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 3.485 1.350 3.745 1.510 ;
        RECT 3.535 1.350 6.095 1.510 ;
        RECT 5.935 0.950 6.095 1.510 ;
        RECT 6.365 4.670 6.625 4.830 ;
        RECT 5.935 4.670 6.575 4.830 ;
        RECT 5.935 1.350 6.575 1.510 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 4.670 6.575 5.830 ;
        RECT 6.415 5.670 12.335 5.830 ;
        RECT 12.125 5.670 12.385 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 7.535 0.450 ;
        RECT 7.375 0.290 7.535 1.110 ;
        RECT 7.375 0.950 8.015 1.110 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 4.495 4.210 8.015 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
        RECT 9.725 0.950 9.985 1.110 ;
        RECT 11.165 1.350 11.425 1.510 ;
        RECT 11.215 1.350 13.295 1.510 ;
        RECT 13.085 1.350 13.345 1.510 ;
        RECT 10.205 0.950 10.465 1.110 ;
        RECT 9.775 0.950 10.415 1.110 ;
  END
END DFQD1
MACRO DFQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_1 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 0.175 0.290 1.775 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 9.245 2.010 9.505 2.170 ;
        RECT 9.295 2.010 9.455 3.610 ;
        RECT 9.245 3.450 9.505 3.610 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 0.335 5.830 ;
        RECT 0.175 5.670 3.695 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.775 3.450 9.935 4.370 ;
        RECT 8.815 4.210 9.935 4.370 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 3.055 2.490 7.535 2.650 ;
        RECT 7.325 2.490 7.585 2.650 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 3.055 2.010 7.535 2.170 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 3.485 4.210 3.745 4.370 ;
        RECT 3.535 4.210 3.695 4.830 ;
        RECT 3.535 4.670 6.095 4.830 ;
        RECT 8.285 0.290 8.545 0.450 ;
        RECT 5.935 0.290 8.495 0.450 ;
        RECT 5.935 0.290 6.095 1.110 ;
        RECT 5.935 4.670 6.095 5.830 ;
        RECT 5.935 5.670 9.455 5.830 ;
        RECT 9.245 5.670 9.505 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 4.495 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 7.855 1.350 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_1
MACRO DFQD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_2 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 1.775 1.110 ;
        RECT 1.615 0.950 1.775 2.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.295 3.450 9.935 3.610 ;
        RECT 9.295 3.450 9.455 4.830 ;
        RECT 8.815 4.670 9.455 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 4.975 0.290 7.535 0.450 ;
        RECT 7.325 0.290 7.585 0.450 ;
        RECT 7.325 4.210 7.585 4.370 ;
        RECT 4.975 4.210 7.535 4.370 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 5.405 1.350 5.665 1.510 ;
        RECT 2.095 1.350 5.615 1.510 ;
        RECT 2.095 0.950 2.255 1.510 ;
        RECT 8.285 2.010 8.545 2.170 ;
        RECT 2.575 2.010 8.495 2.170 ;
        RECT 2.575 2.010 2.735 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 5.455 1.350 5.615 2.170 ;
        RECT 8.335 2.010 8.495 5.830 ;
        RECT 8.335 5.670 9.455 5.830 ;
        RECT 9.245 5.670 9.505 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 3.535 5.670 8.495 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 6.365 3.450 6.625 3.610 ;
        RECT 6.415 3.450 8.015 3.610 ;
        RECT 7.855 3.450 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_2
MACRO DFQD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_3 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 2.970 1.345 3.130 ;
        RECT 1.135 2.970 1.295 3.610 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.950 12.865 1.110 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 12.655 0.950 12.815 4.830 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 14.280 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 14.280 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 9.245 0.290 9.505 0.450 ;
        RECT 4.015 0.290 9.455 0.450 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 2.575 0.950 4.175 1.110 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 1.775 2.170 ;
        RECT 1.615 2.010 1.775 4.830 ;
        RECT 1.615 4.670 2.255 4.830 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 0.655 2.490 2.255 2.650 ;
        RECT 0.605 2.490 0.865 2.650 ;
        RECT 8.765 0.950 9.025 1.110 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 8.815 0.950 11.375 1.110 ;
        RECT 11.215 0.290 11.375 1.110 ;
        RECT 11.165 0.290 11.425 0.450 ;
        RECT 9.775 0.950 9.935 3.610 ;
        RECT 9.775 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
        RECT 9.295 3.450 9.935 3.610 ;
        RECT 9.295 3.450 9.455 4.830 ;
        RECT 8.815 4.670 9.455 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
        RECT 7.325 2.010 7.585 2.170 ;
        RECT 4.975 2.010 7.535 2.170 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.175 0.290 3.695 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 8.495 5.170 ;
        RECT 8.335 3.450 8.495 5.170 ;
        RECT 8.285 3.450 8.545 3.610 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 3.535 5.010 3.695 5.830 ;
        RECT 7.805 0.950 8.065 1.110 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 6.365 1.350 6.625 1.510 ;
        RECT 6.415 1.350 8.015 1.510 ;
        RECT 7.855 0.950 8.015 1.510 ;
        RECT 7.855 1.350 8.015 4.830 ;
        RECT 11.645 0.950 11.905 1.110 ;
        RECT 10.205 1.350 10.465 1.510 ;
        RECT 10.255 1.350 12.335 1.510 ;
        RECT 12.175 0.290 12.335 1.510 ;
        RECT 12.175 0.290 13.295 0.450 ;
        RECT 13.085 0.290 13.345 0.450 ;
        RECT 11.695 0.950 11.855 1.510 ;
  END
END DFQD1_3
#--------EOF---------

MACRO FILL1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL1 0 0 ; 
  SIZE 0.340 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 0.340 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 0.340 0.100 ;
    END 
  END vss 
END FILL1
#--------EOF---------

MACRO FILL1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL1 0 0 ; 
  SIZE 0.340 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 0.340 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 0.340 0.100 ;
    END 
  END vss 
END FILL1
#--------EOF---------

MACRO FILL2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL2 0 0 ; 
  SIZE 0.680 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 0.680 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 0.680 0.100 ;
    END 
  END vss 
END FILL2
#--------EOF---------

MACRO FILL2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL2 0 0 ; 
  SIZE 0.680 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 0.680 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 0.680 0.100 ;
    END 
  END vss 
END FILL2
#--------EOF---------

MACRO FILL4
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL4 0 0 ; 
  SIZE 1.360 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 1.360 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 1.360 0.100 ;
    END 
  END vss 
END FILL4
#--------EOF---------

MACRO FILL4
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL4 0 0 ; 
  SIZE 1.360 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 1.360 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 1.360 0.100 ;
    END 
  END vss 
END FILL4
#--------EOF---------

MACRO FILL8
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL8 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END FILL8
#--------EOF---------

MACRO FILL8
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL8 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END FILL8
#--------EOF---------

MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1
MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1
MACRO INVD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_1
MACRO INVD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_2 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_2
MACRO INVD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_3 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_3
#--------EOF---------

MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1
MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1
MACRO INVD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_1
MACRO INVD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_2 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_2
MACRO INVD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_3 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
END INVD1_3
#--------EOF---------

MACRO MUX2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 1.350 2.735 2.170 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 1.350 1.775 2.170 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 0.655 0.290 4.655 0.450 ;
        RECT 4.495 0.290 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 5.405 2.010 5.665 2.170 ;
        RECT 5.455 2.010 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 2.170 ;
        RECT 1.085 2.010 1.345 2.170 ;
        RECT 1.085 3.450 1.345 3.610 ;
        RECT 1.135 3.450 1.295 4.830 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.015 0.950 4.175 3.610 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 0.175 2.490 2.735 2.650 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 4.015 2.490 4.175 5.170 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.925 0.290 5.185 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 3.005 5.670 3.265 5.830 ;
        RECT 3.055 5.670 5.135 5.830 ;
        RECT 4.975 5.010 5.135 5.830 ;
  END
END MUX2D1
MACRO MUX2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 3.055 2.970 4.655 3.130 ;
        RECT 3.005 2.970 3.265 3.130 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 2.095 5.010 4.655 5.170 ;
        RECT 4.495 4.210 4.655 5.170 ;
        RECT 4.495 4.210 5.135 4.370 ;
        RECT 4.925 4.210 5.185 4.370 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.650 ;
        RECT 2.575 2.490 3.215 2.650 ;
        RECT 2.575 2.490 2.735 4.830 ;
        RECT 2.575 4.670 3.215 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 1.615 2.010 2.735 2.170 ;
        RECT 1.615 2.010 1.775 3.610 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 4.975 0.950 5.615 1.110 ;
        RECT 5.455 0.950 5.615 5.170 ;
        RECT 4.975 5.010 5.615 5.170 ;
        RECT 1.565 5.670 1.825 5.830 ;
        RECT 1.615 5.670 5.135 5.830 ;
        RECT 4.975 5.010 5.135 5.830 ;
  END
END MUX2D1_1
MACRO MUX2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.935 0.070 6.095 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 3.215 4.830 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 4.015 0.290 5.135 0.450 ;
        RECT 4.925 0.290 5.185 0.450 ;
        RECT 4.015 0.950 4.175 5.170 ;
        RECT 0.655 2.970 4.175 3.130 ;
        RECT 0.655 2.970 0.815 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
        RECT 0.175 0.950 0.335 3.130 ;
        RECT 0.175 2.970 0.815 3.130 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 2.170 ;
        RECT 1.085 2.010 1.345 2.170 ;
        RECT 1.085 3.450 1.345 3.610 ;
        RECT 1.135 3.450 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.445 0.950 4.705 1.110 ;
        RECT 4.495 0.950 5.135 1.110 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 3.535 0.290 3.695 2.650 ;
        RECT 3.485 2.490 3.745 2.650 ;
        RECT 4.975 0.950 5.135 5.170 ;
  END
END MUX2D1_2
MACRO MUX2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 2.735 1.110 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 5.010 4.175 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 3.215 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 5.170 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 2.095 2.970 4.655 3.130 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 2.525 4.210 2.785 4.370 ;
        RECT 2.575 4.210 2.735 5.170 ;
        RECT 2.575 5.010 3.695 5.170 ;
        RECT 3.535 4.670 3.695 5.170 ;
        RECT 3.535 4.670 5.135 4.830 ;
        RECT 4.975 4.670 5.135 5.170 ;
        RECT 4.975 0.950 5.135 4.830 ;
  END
END MUX2D1_3
#--------EOF---------

MACRO MUX2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 1.350 2.735 2.170 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 1.350 1.775 2.170 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 0.655 0.290 4.655 0.450 ;
        RECT 4.495 0.290 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 5.405 2.010 5.665 2.170 ;
        RECT 5.455 2.010 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 2.170 ;
        RECT 1.085 2.010 1.345 2.170 ;
        RECT 1.085 3.450 1.345 3.610 ;
        RECT 1.135 3.450 1.295 4.830 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.015 0.950 4.175 3.610 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 0.175 2.490 2.735 2.650 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 4.015 2.490 4.175 5.170 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.925 0.290 5.185 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 3.005 5.670 3.265 5.830 ;
        RECT 3.055 5.670 5.135 5.830 ;
        RECT 4.975 5.010 5.135 5.830 ;
  END
END MUX2D1
MACRO MUX2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 3.055 2.970 4.655 3.130 ;
        RECT 3.005 2.970 3.265 3.130 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 2.095 5.010 4.655 5.170 ;
        RECT 4.495 4.210 4.655 5.170 ;
        RECT 4.495 4.210 5.135 4.370 ;
        RECT 4.925 4.210 5.185 4.370 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.650 ;
        RECT 2.575 2.490 3.215 2.650 ;
        RECT 2.575 2.490 2.735 4.830 ;
        RECT 2.575 4.670 3.215 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 1.615 2.010 2.735 2.170 ;
        RECT 1.615 2.010 1.775 3.610 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 4.975 0.950 5.615 1.110 ;
        RECT 5.455 0.950 5.615 5.170 ;
        RECT 4.975 5.010 5.615 5.170 ;
        RECT 1.565 5.670 1.825 5.830 ;
        RECT 1.615 5.670 5.135 5.830 ;
        RECT 4.975 5.010 5.135 5.830 ;
  END
END MUX2D1_1
MACRO MUX2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.935 0.070 6.095 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 3.215 4.830 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 4.015 0.290 5.135 0.450 ;
        RECT 4.925 0.290 5.185 0.450 ;
        RECT 4.015 0.950 4.175 5.170 ;
        RECT 0.655 2.970 4.175 3.130 ;
        RECT 0.655 2.970 0.815 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
        RECT 0.175 0.950 0.335 3.130 ;
        RECT 0.175 2.970 0.815 3.130 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 2.170 ;
        RECT 1.085 2.010 1.345 2.170 ;
        RECT 1.085 3.450 1.345 3.610 ;
        RECT 1.135 3.450 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.445 0.950 4.705 1.110 ;
        RECT 4.495 0.950 5.135 1.110 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 3.535 0.290 3.695 2.650 ;
        RECT 3.485 2.490 3.745 2.650 ;
        RECT 4.975 0.950 5.135 5.170 ;
  END
END MUX2D1_2
MACRO MUX2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 2.735 1.110 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 5.010 4.175 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 3.215 4.830 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 5.170 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 2.095 2.970 4.655 3.130 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 2.525 4.210 2.785 4.370 ;
        RECT 2.575 4.210 2.735 5.170 ;
        RECT 2.575 5.010 3.695 5.170 ;
        RECT 3.535 4.670 3.695 5.170 ;
        RECT 3.535 4.670 5.135 4.830 ;
        RECT 4.975 4.670 5.135 5.170 ;
        RECT 4.975 0.950 5.135 4.830 ;
  END
END MUX2D1_3
#--------EOF---------

MACRO ND2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 1.135 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1
MACRO ND2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_1
MACRO ND2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_2
MACRO ND2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_3
#--------EOF---------

MACRO ND2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 1.135 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1
MACRO ND2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_1
MACRO ND2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_2
MACRO ND2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END ND2D1_3
#--------EOF---------

MACRO ND3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END ND3D1
MACRO ND3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_1 0 0 ; 
  SIZE 3.400 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.400 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.400 0.100 ;
    END 
  END vss 
END ND3D1_1
MACRO ND3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_2 0 0 ; 
  SIZE 4.760 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.760 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.760 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 0.175 0.290 4.175 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END ND3D1_2
MACRO ND3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END ND3D1_3
#--------EOF---------

MACRO ND3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END ND3D1
MACRO ND3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_1 0 0 ; 
  SIZE 3.400 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.400 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.400 0.100 ;
    END 
  END vss 
END ND3D1_1
MACRO ND3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_2 0 0 ; 
  SIZE 4.760 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.760 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.760 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 0.175 0.290 4.175 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END ND3D1_2
MACRO ND3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END ND3D1_3
#--------EOF---------

MACRO ND4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 0.950 3.215 4.370 ;
        RECT 3.055 4.210 4.175 4.370 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 0.175 0.290 4.175 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END ND4D1
MACRO ND4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
        RECT 1.135 4.210 4.175 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.535 4.670 4.175 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 5.135 6.050 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 5.135 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
  END
END ND4D1_1
MACRO ND4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
END ND4D1_2
MACRO ND4D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 4.975 0.950 5.135 4.370 ;
        RECT 4.015 4.210 5.135 4.370 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 1.135 4.210 4.175 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 5.135 6.050 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 3.215 1.110 ;
  END
END ND4D1_3
#--------EOF---------

MACRO ND4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.055 0.950 3.215 4.370 ;
        RECT 3.055 4.210 4.175 4.370 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 1.135 4.210 3.215 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 0.175 0.290 4.175 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END ND4D1
MACRO ND4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
        RECT 1.135 4.210 4.175 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.535 4.670 4.175 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 5.135 6.050 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 0.175 0.290 5.135 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
  END
END ND4D1_1
MACRO ND4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
END ND4D1_2
MACRO ND4D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 4.975 0.950 5.135 4.370 ;
        RECT 4.015 4.210 5.135 4.370 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 1.135 4.210 4.175 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 5.135 6.050 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 3.215 1.110 ;
  END
END ND4D1_3
#--------EOF---------

MACRO NR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 0.175 4.670 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1
MACRO NR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_1
MACRO NR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_2
MACRO NR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_3
#--------EOF---------

MACRO NR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 0.175 4.670 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 4.670 2.255 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1
MACRO NR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.095 0.070 2.255 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_1
MACRO NR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_2
MACRO NR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 2.720 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 2.720 0.100 ;
    END 
  END vss 
END NR2D1_3
#--------EOF---------

MACRO NR3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 1.615 0.290 1.775 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 2.735 1.110 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 3.055 0.950 3.215 3.610 ;
        RECT 1.135 3.450 3.215 3.610 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 0.175 5.010 8.015 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
  END
END NR3D1
MACRO NR3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_1 0 0 ; 
  SIZE 10.540 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 1.350 3.695 2.170 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 5.615 2.650 ;
        RECT 5.405 2.490 5.665 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 10.540 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 10.540 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 8.815 4.670 8.975 5.170 ;
        RECT 2.095 5.010 8.975 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 9.775 4.210 9.935 4.830 ;
        RECT 6.895 4.210 9.935 4.370 ;
        RECT 6.895 4.210 7.055 4.830 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 4.670 5.135 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
        RECT 1.615 4.210 3.215 4.370 ;
        RECT 1.615 4.210 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR3D1_1
MACRO NR3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_2 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 0.335 4.370 ;
        RECT 0.175 4.210 1.295 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 0.175 5.010 8.015 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
  END
END NR3D1_2
MACRO NR3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_3 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 1.135 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 3.055 5.010 8.015 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 2.575 4.210 4.175 4.370 ;
        RECT 2.575 4.210 2.735 5.170 ;
        RECT 0.175 5.010 2.735 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR3D1_3
#--------EOF---------

MACRO NR3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 1.615 0.290 1.775 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 2.735 1.110 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 3.055 0.950 3.215 3.610 ;
        RECT 1.135 3.450 3.215 3.610 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 0.175 5.010 8.015 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
  END
END NR3D1
MACRO NR3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_1 0 0 ; 
  SIZE 10.540 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 1.350 3.695 2.170 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 5.615 2.650 ;
        RECT 5.405 2.490 5.665 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 0.950 3.215 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 10.540 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 10.540 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 8.815 4.670 8.975 5.170 ;
        RECT 2.095 5.010 8.975 5.170 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 9.775 4.210 9.935 4.830 ;
        RECT 6.895 4.210 9.935 4.370 ;
        RECT 6.895 4.210 7.055 4.830 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 4.670 5.135 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.055 4.210 3.215 4.830 ;
        RECT 1.615 4.210 3.215 4.370 ;
        RECT 1.615 4.210 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR3D1_1
MACRO NR3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_2 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 0.175 0.950 0.335 4.370 ;
        RECT 0.175 4.210 1.295 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 0.175 5.010 8.015 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 4.175 4.830 ;
  END
END NR3D1_2
MACRO NR3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_3 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 3.215 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 1.135 0.950 2.255 1.110 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 9.520 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 9.520 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 7.855 4.670 8.015 5.170 ;
        RECT 3.055 5.010 8.015 5.170 ;
        RECT 3.055 4.670 3.215 5.170 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 8.815 4.210 8.975 4.830 ;
        RECT 5.935 4.210 8.975 4.370 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 2.575 4.210 4.175 4.370 ;
        RECT 2.575 4.210 2.735 5.170 ;
        RECT 0.175 5.010 2.735 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR3D1_3
#--------EOF---------

MACRO NR4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 0.655 0.290 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 4.015 3.450 6.575 3.610 ;
        RECT 6.365 3.450 6.625 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.450 8.065 3.610 ;
        RECT 7.855 3.450 12.335 3.610 ;
        RECT 12.125 3.450 12.385 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 13.260 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 13.260 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 4.670 11.855 4.830 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 12.175 4.670 12.815 4.830 ;
        RECT 12.175 4.210 12.335 4.830 ;
        RECT 7.855 4.210 12.335 4.370 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.615 4.670 3.215 4.830 ;
        RECT 1.615 4.670 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 4.975 4.670 6.575 4.830 ;
        RECT 6.415 4.210 6.575 4.830 ;
        RECT 6.415 4.210 7.535 4.370 ;
        RECT 7.325 4.210 7.585 4.370 ;
        RECT 7.325 5.010 7.585 5.170 ;
        RECT 7.375 5.010 9.935 5.170 ;
        RECT 9.775 4.670 9.935 5.170 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 2.095 4.210 6.095 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END NR4D1
MACRO NR4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_1 0 0 ; 
  SIZE 12.240 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 5.615 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 3.450 7.105 3.610 ;
        RECT 6.895 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 3.215 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 12.240 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 12.240 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 10.685 4.670 10.945 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 4.670 10.895 4.830 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 11.215 4.670 11.855 4.830 ;
        RECT 11.215 4.210 11.375 4.830 ;
        RECT 6.895 4.210 11.375 4.370 ;
        RECT 6.895 4.210 7.055 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 4.015 4.670 5.615 4.830 ;
        RECT 5.455 4.210 5.615 4.830 ;
        RECT 5.455 4.210 6.575 4.370 ;
        RECT 6.365 4.210 6.625 4.370 ;
        RECT 6.365 5.010 6.625 5.170 ;
        RECT 6.415 5.010 8.975 5.170 ;
        RECT 8.815 4.670 8.975 5.170 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 1.615 4.210 5.135 4.370 ;
        RECT 1.615 4.210 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR4D1_1
MACRO NR4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_2 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 4.655 5.830 ;
        RECT 3.535 5.670 4.655 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 4.445 5.670 4.705 5.830 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.655 0.290 3.695 0.450 ;
        RECT 0.655 0.290 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 3.695 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.450 8.065 3.610 ;
        RECT 7.855 3.450 12.335 3.610 ;
        RECT 12.125 3.450 12.385 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 13.260 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 13.260 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 4.670 11.855 4.830 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 12.175 4.670 12.815 4.830 ;
        RECT 12.175 4.210 12.335 4.830 ;
        RECT 7.855 4.210 12.335 4.370 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.175 4.670 3.215 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 2.095 4.210 2.735 4.370 ;
        RECT 2.525 4.210 2.785 4.370 ;
        RECT 7.325 5.010 7.585 5.170 ;
        RECT 7.375 5.010 9.935 5.170 ;
        RECT 9.775 4.670 9.935 5.170 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 6.095 4.830 ;
  END
END NR4D1_2
#--------EOF---------

MACRO NR4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 0.655 0.290 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 4.015 3.450 6.575 3.610 ;
        RECT 6.365 3.450 6.625 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.450 8.065 3.610 ;
        RECT 7.855 3.450 12.335 3.610 ;
        RECT 12.125 3.450 12.385 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 13.260 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 13.260 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 4.670 11.855 4.830 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 12.175 4.670 12.815 4.830 ;
        RECT 12.175 4.210 12.335 4.830 ;
        RECT 7.855 4.210 12.335 4.370 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 1.615 4.670 3.215 4.830 ;
        RECT 1.615 4.670 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 4.975 4.670 6.575 4.830 ;
        RECT 6.415 4.210 6.575 4.830 ;
        RECT 6.415 4.210 7.535 4.370 ;
        RECT 7.325 4.210 7.585 4.370 ;
        RECT 7.325 5.010 7.585 5.170 ;
        RECT 7.375 5.010 9.935 5.170 ;
        RECT 9.775 4.670 9.935 5.170 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 5.935 4.210 6.095 4.830 ;
        RECT 2.095 4.210 6.095 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END NR4D1
MACRO NR4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_1 0 0 ; 
  SIZE 12.240 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 3.450 3.265 3.610 ;
        RECT 3.055 3.450 5.615 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 3.450 7.105 3.610 ;
        RECT 6.895 3.450 11.375 3.610 ;
        RECT 11.165 3.450 11.425 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 3.215 1.110 ;
        RECT 1.135 0.950 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 12.240 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 12.240 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 10.685 4.670 10.945 4.830 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 4.670 10.895 4.830 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 11.215 4.670 11.855 4.830 ;
        RECT 11.215 4.210 11.375 4.830 ;
        RECT 6.895 4.210 11.375 4.370 ;
        RECT 6.895 4.210 7.055 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 8.765 4.670 9.025 4.830 ;
        RECT 4.015 4.670 5.615 4.830 ;
        RECT 5.455 4.210 5.615 4.830 ;
        RECT 5.455 4.210 6.575 4.370 ;
        RECT 6.365 4.210 6.625 4.370 ;
        RECT 6.365 5.010 6.625 5.170 ;
        RECT 6.415 5.010 8.975 5.170 ;
        RECT 8.815 4.670 8.975 5.170 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 4.975 4.210 5.135 4.830 ;
        RECT 1.615 4.210 5.135 4.370 ;
        RECT 1.615 4.210 1.775 5.170 ;
        RECT 0.175 5.010 1.775 5.170 ;
        RECT 0.175 4.670 0.335 5.170 ;
  END
END NR4D1_1
MACRO NR4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_2 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 4.655 5.830 ;
        RECT 3.535 5.670 4.655 5.830 ;
        RECT 3.485 5.670 3.745 5.830 ;
        RECT 4.445 5.670 4.705 5.830 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.655 0.290 3.695 0.450 ;
        RECT 0.655 0.290 0.815 3.610 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 3.695 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.450 8.065 3.610 ;
        RECT 7.855 3.450 12.335 3.610 ;
        RECT 12.125 3.450 12.385 3.610 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 1.135 0.950 4.175 1.110 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 13.260 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 13.260 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.670 11.905 4.830 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 4.670 11.855 4.830 ;
        RECT 12.605 4.670 12.865 4.830 ;
        RECT 7.805 4.670 8.065 4.830 ;
        RECT 12.175 4.670 12.815 4.830 ;
        RECT 12.175 4.210 12.335 4.830 ;
        RECT 7.855 4.210 12.335 4.370 ;
        RECT 7.855 4.210 8.015 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.175 4.670 3.215 4.830 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 9.725 4.670 9.985 4.830 ;
        RECT 2.095 4.210 2.255 4.830 ;
        RECT 2.095 4.210 2.735 4.370 ;
        RECT 2.525 4.210 2.785 4.370 ;
        RECT 7.325 5.010 7.585 5.170 ;
        RECT 7.375 5.010 9.935 5.170 ;
        RECT 9.775 4.670 9.935 5.170 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 4.670 6.095 4.830 ;
  END
END NR4D1_2
#--------EOF---------

MACRO OA21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.535 0.950 4.175 1.110 ;
        RECT 3.485 0.950 3.745 1.110 ;
        RECT 0.175 0.950 0.335 4.370 ;
        RECT 0.175 4.210 1.295 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 1.135 0.290 5.135 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 4.175 5.170 ;
        RECT 4.015 4.670 4.175 5.170 ;
  END
END OA21D1
MACRO OA21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 2.575 2.490 2.735 3.130 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 2.095 2.010 3.215 2.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
  END
END OA21D1_1
MACRO OA21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 2.650 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 4.015 3.450 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 0.655 2.970 4.655 3.130 ;
        RECT 0.655 2.970 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 1.135 2.970 1.775 3.130 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 0.175 0.290 2.255 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END OA21D1_2
MACRO OA21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 3.485 4.670 3.745 4.830 ;
        RECT 3.055 4.670 3.695 4.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OA21D1_3
#--------EOF---------

MACRO OA21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.010 4.705 2.170 ;
        RECT 4.495 2.010 4.655 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 3.535 0.950 4.175 1.110 ;
        RECT 3.485 0.950 3.745 1.110 ;
        RECT 0.175 0.950 0.335 4.370 ;
        RECT 0.175 4.210 1.295 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 1.135 0.290 5.135 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 0.175 4.670 0.335 5.170 ;
        RECT 0.175 5.010 4.175 5.170 ;
        RECT 4.015 4.670 4.175 5.170 ;
  END
END OA21D1
MACRO OA21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.490 2.785 2.650 ;
        RECT 2.575 2.490 2.735 3.130 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 2.095 2.010 3.215 2.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 1.135 0.290 1.295 1.110 ;
  END
END OA21D1_1
MACRO OA21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 2.650 ;
        RECT 3.965 2.490 4.225 2.650 ;
        RECT 3.965 3.450 4.225 3.610 ;
        RECT 4.015 3.450 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 4.670 3.215 4.830 ;
        RECT 4.445 2.970 4.705 3.130 ;
        RECT 0.655 2.970 4.655 3.130 ;
        RECT 0.655 2.970 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 1.135 2.970 1.775 3.130 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 0.175 0.290 2.255 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END OA21D1_2
MACRO OA21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 4.670 4.225 4.830 ;
        RECT 4.015 0.950 4.175 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 5.440 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 5.440 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 3.485 4.670 3.745 4.830 ;
        RECT 3.055 4.670 3.695 4.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OA21D1_3
#--------EOF---------

MACRO OAI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1
MACRO OAI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 0.175 0.290 2.255 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END OAI21D1_1
MACRO OAI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 3.215 4.830 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.525 4.670 2.785 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1_2
MACRO OAI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 0.175 0.950 0.335 1.510 ;
        RECT 0.175 1.350 2.255 1.510 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1_3
#--------EOF---------

MACRO OAI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 2.095 0.950 2.255 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 1.135 4.210 1.295 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.070 0.335 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1
MACRO OAI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 4.670 3.215 6.050 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.175 4.670 0.335 6.050 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.055 0.070 3.215 1.110 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 0.175 0.290 2.255 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
  END
END OAI21D1_1
MACRO OAI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 0.175 0.950 0.335 4.830 ;
        RECT 0.175 4.670 3.215 4.830 ;
        RECT 2.095 0.950 2.735 1.110 ;
        RECT 2.525 0.950 2.785 1.110 ;
        RECT 2.525 4.670 2.785 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1_2
MACRO OAI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 2.650 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 0.175 0.950 0.335 1.510 ;
        RECT 0.175 1.350 2.255 1.510 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.135 0.290 3.215 0.450 ;
        RECT 3.055 0.290 3.215 1.110 ;
  END
END OAI21D1_3
#--------EOF---------

MACRO OR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 0.175 2.970 2.735 3.130 ;
        RECT 0.175 2.970 0.335 4.830 ;
        RECT 1.135 0.950 1.295 3.130 ;
  END
END OR2D1
MACRO OR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.525 4.670 2.785 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END OR2D1_1
MACRO OR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 0.290 2.305 0.450 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
  END
END OR2D1_2
MACRO OR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.175 0.290 3.695 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 2.095 0.290 2.255 4.830 ;
        RECT 2.095 0.290 2.255 1.110 ;
  END
END OR2D1_3
#--------EOF---------

MACRO OR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 3.740 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 3.740 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 0.175 2.970 2.735 3.130 ;
        RECT 0.175 2.970 0.335 4.830 ;
        RECT 1.135 0.950 1.295 3.130 ;
  END
END OR2D1
MACRO OR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.525 4.670 2.785 4.830 ;
        RECT 2.095 4.670 2.735 4.830 ;
        RECT 1.135 0.950 1.295 4.370 ;
        RECT 1.135 4.210 2.255 4.370 ;
        RECT 2.095 4.210 2.255 4.830 ;
  END
END OR2D1_1
MACRO OR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 2.045 0.290 2.305 0.450 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.950 2.255 4.830 ;
        RECT 0.175 4.670 2.255 4.830 ;
        RECT 0.175 0.950 2.255 1.110 ;
  END
END OR2D1_2
MACRO OR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 1.775 2.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 4.670 3.265 4.830 ;
        RECT 3.055 0.950 3.215 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 4.420 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 4.420 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 0.175 0.290 3.695 0.450 ;
        RECT 0.175 0.290 0.335 1.110 ;
        RECT 2.095 0.290 2.255 4.830 ;
        RECT 2.095 0.290 2.255 1.110 ;
  END
END OR2D1_3
#--------EOF---------

MACRO TAPCELL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL 0 0 ; 
  SIZE 2.380 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 4.750 0.600 4.910 ;
        RECT 0.390 4.750 0.550 6.050 ;
        RECT 0.820 4.750 1.080 4.910 ;
        RECT 0.870 4.750 1.030 6.050 ;
        RECT 1.300 4.750 1.560 4.910 ;
        RECT 1.350 4.750 1.510 6.050 ;
        RECT 0.000 6.020 2.380 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 0.870 0.600 1.030 ;
        RECT 0.390 0.070 0.550 1.030 ;
        RECT 0.820 0.870 1.080 1.030 ;
        RECT 0.870 0.070 1.030 1.030 ;
        RECT 1.300 0.870 1.560 1.030 ;
        RECT 1.350 0.070 1.510 1.030 ;
        RECT 0.000 -0.100 2.380 0.100 ;
    END 
  END vss 
END TAPCELL
#--------EOF---------

MACRO TAPCELL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL 0 0 ; 
  SIZE 2.380 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 4.750 0.600 4.910 ;
        RECT 0.390 4.750 0.550 6.050 ;
        RECT 0.820 4.750 1.080 4.910 ;
        RECT 0.870 4.750 1.030 6.050 ;
        RECT 1.300 4.750 1.560 4.910 ;
        RECT 1.350 4.750 1.510 6.050 ;
        RECT 0.000 6.020 2.380 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 0.870 0.600 1.030 ;
        RECT 0.390 0.070 0.550 1.030 ;
        RECT 0.820 0.870 1.080 1.030 ;
        RECT 0.870 0.070 1.030 1.030 ;
        RECT 1.300 0.870 1.560 1.030 ;
        RECT 1.350 0.070 1.510 1.030 ;
        RECT 0.000 -0.100 2.380 0.100 ;
    END 
  END vss 
END TAPCELL
#--------EOF---------

MACRO TIEH
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEH 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 0.655 4.670 0.815 5.170 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 0.815 1.110 ;
        RECT 0.655 0.290 0.815 1.110 ;
        RECT 0.605 0.290 0.865 0.450 ;
  END
END TIEH
#--------EOF---------

MACRO TIEH
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEH 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 4.670 0.815 4.830 ;
        RECT 0.655 4.670 0.815 5.170 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 0.175 0.950 0.815 1.110 ;
        RECT 0.655 0.290 0.815 1.110 ;
        RECT 0.605 0.290 0.865 0.450 ;
  END
END TIEH
#--------EOF---------

MACRO TIEL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEL 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 0.950 0.815 1.110 ;
        RECT 0.655 0.950 0.815 1.510 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
  END
END TIEL
#--------EOF---------

MACRO TIEL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEL 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 0.950 0.815 1.110 ;
        RECT 0.655 0.950 0.815 1.510 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 4.670 1.295 6.050 ;
        RECT 0.000 6.020 1.700 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.135 0.070 1.295 1.110 ;
        RECT 0.000 -0.100 1.700 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.670 0.385 4.830 ;
        RECT 0.605 3.450 0.865 3.610 ;
        RECT 0.655 3.450 0.815 4.830 ;
        RECT 0.175 4.670 0.815 4.830 ;
  END
END TIEL
#--------EOF---------

MACRO XNR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 4.655 1.110 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 5.010 1.295 5.830 ;
        RECT 1.085 5.670 1.345 5.830 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 4.210 3.265 4.370 ;
        RECT 3.055 4.210 3.215 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 2.095 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 2.095 5.010 2.255 5.830 ;
        RECT 2.095 5.670 6.575 5.830 ;
        RECT 6.365 5.670 6.625 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.975 0.950 5.135 3.130 ;
        RECT 1.615 2.970 5.135 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 4.975 2.970 5.135 5.170 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 2.575 2.970 5.135 3.130 ;
  END
END XNR2D1
MACRO XNR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 5.010 4.175 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 0.655 0.290 3.215 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 3.055 5.010 3.215 5.830 ;
        RECT 0.655 5.670 3.215 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 3.005 2.970 3.265 3.130 ;
        RECT 3.055 2.970 3.215 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 2.095 2.490 3.215 2.650 ;
        RECT 3.055 2.490 3.215 3.130 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.975 0.950 5.135 1.510 ;
        RECT 2.575 1.350 5.135 1.510 ;
        RECT 2.575 1.350 2.735 2.170 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 4.975 1.350 5.135 5.170 ;
  END
END XNR2D1_1
MACRO XNR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 1.615 2.970 3.215 3.130 ;
        RECT 3.005 2.970 3.265 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 3.215 2.170 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 5.615 0.450 ;
        RECT 5.405 0.290 5.665 0.450 ;
        RECT 5.455 0.290 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
        RECT 2.095 4.670 4.175 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 3.965 4.210 4.225 4.370 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.975 5.010 5.135 5.830 ;
        RECT 0.175 5.670 5.135 5.830 ;
        RECT 0.175 5.010 0.335 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 3.485 2.490 3.745 2.650 ;
        RECT 1.135 2.490 3.695 2.650 ;
        RECT 1.135 2.490 1.295 5.170 ;
        RECT 1.135 0.950 1.295 2.650 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 0.950 4.175 1.510 ;
        RECT 1.615 1.350 4.175 1.510 ;
        RECT 1.615 0.290 1.775 1.510 ;
        RECT 0.655 0.290 1.775 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 2.095 1.350 2.255 2.170 ;
        RECT 2.045 2.010 2.305 2.170 ;
        RECT 4.015 1.350 4.655 1.510 ;
        RECT 4.495 1.350 4.655 5.170 ;
        RECT 4.015 5.010 4.655 5.170 ;
  END
END XNR2D1_2
MACRO XNR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 1.615 0.290 3.695 0.450 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 3.485 4.210 3.745 4.370 ;
        RECT 0.655 4.210 3.695 4.370 ;
        RECT 0.605 4.210 0.865 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 4.655 1.110 ;
        RECT 4.495 0.290 4.655 1.110 ;
        RECT 4.495 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 4.015 0.950 4.175 4.830 ;
        RECT 2.095 4.670 4.175 4.830 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 6.845 5.010 7.105 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 5.455 0.950 7.055 1.110 ;
        RECT 5.455 0.950 5.615 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 4.445 5.010 4.705 5.170 ;
        RECT 0.175 5.010 4.655 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.495 5.010 7.055 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
  END
END XNR2D1_3
#--------EOF---------

MACRO XNR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.290 4.705 0.450 ;
        RECT 4.495 0.290 4.655 1.110 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 5.010 1.295 5.830 ;
        RECT 1.085 5.670 1.345 5.830 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.950 3.215 2.170 ;
        RECT 3.005 2.010 3.265 2.170 ;
        RECT 3.005 4.210 3.265 4.370 ;
        RECT 3.055 4.210 3.215 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 2.095 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 2.095 5.010 2.255 5.830 ;
        RECT 2.095 5.670 6.575 5.830 ;
        RECT 6.365 5.670 6.625 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.975 0.950 5.135 3.130 ;
        RECT 1.615 2.970 5.135 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 4.975 2.970 5.135 5.170 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 2.575 2.970 5.135 3.130 ;
  END
END XNR2D1
MACRO XNR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.495 2.490 4.655 4.370 ;
        RECT 4.445 4.210 4.705 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.010 3.745 2.170 ;
        RECT 3.535 2.010 3.695 3.610 ;
        RECT 3.485 3.450 3.745 3.610 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 5.010 4.175 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 4.015 0.070 4.175 1.110 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.290 3.215 1.110 ;
        RECT 0.655 0.290 3.215 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 3.055 5.010 3.215 5.830 ;
        RECT 0.655 5.670 3.215 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 3.005 2.970 3.265 3.130 ;
        RECT 3.055 2.970 3.215 4.830 ;
        RECT 2.095 4.670 3.215 4.830 ;
        RECT 2.095 4.670 2.255 5.170 ;
        RECT 2.095 0.950 2.255 2.650 ;
        RECT 2.095 2.490 3.215 2.650 ;
        RECT 3.055 2.490 3.215 3.130 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 4.975 0.950 5.135 1.510 ;
        RECT 2.575 1.350 5.135 1.510 ;
        RECT 2.575 1.350 2.735 2.170 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 4.975 1.350 5.135 5.170 ;
  END
END XNR2D1_1
MACRO XNR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 1.615 2.970 3.215 3.130 ;
        RECT 3.005 2.970 3.265 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 3.215 2.170 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 5.010 6.145 5.170 ;
        RECT 5.935 5.010 6.095 6.050 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 5.615 0.450 ;
        RECT 5.405 0.290 5.665 0.450 ;
        RECT 5.455 0.290 5.615 4.370 ;
        RECT 5.405 4.210 5.665 4.370 ;
        RECT 2.095 4.670 4.175 4.830 ;
        RECT 4.015 4.210 4.175 4.830 ;
        RECT 3.965 4.210 4.225 4.370 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.975 5.010 5.135 5.830 ;
        RECT 0.175 5.670 5.135 5.830 ;
        RECT 0.175 5.010 0.335 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 3.485 2.490 3.745 2.650 ;
        RECT 1.135 2.490 3.695 2.650 ;
        RECT 1.135 2.490 1.295 5.170 ;
        RECT 1.135 0.950 1.295 2.650 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 4.015 0.950 4.175 1.510 ;
        RECT 1.615 1.350 4.175 1.510 ;
        RECT 1.615 0.290 1.775 1.510 ;
        RECT 0.655 0.290 1.775 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 2.095 1.350 2.255 2.170 ;
        RECT 2.045 2.010 2.305 2.170 ;
        RECT 4.015 1.350 4.655 1.510 ;
        RECT 4.495 1.350 4.655 5.170 ;
        RECT 4.015 5.010 4.655 5.170 ;
  END
END XNR2D1_2
MACRO XNR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.290 3.745 0.450 ;
        RECT 1.615 0.290 3.695 0.450 ;
        RECT 1.565 0.290 1.825 0.450 ;
        RECT 3.485 4.210 3.745 4.370 ;
        RECT 0.655 4.210 3.695 4.370 ;
        RECT 0.605 4.210 0.865 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 4.670 2.305 4.830 ;
        RECT 2.095 0.950 4.655 1.110 ;
        RECT 4.495 0.290 4.655 1.110 ;
        RECT 4.495 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 4.015 0.950 4.175 4.830 ;
        RECT 2.095 4.670 4.175 4.830 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 6.845 5.010 7.105 5.170 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 5.455 0.950 7.055 1.110 ;
        RECT 5.455 0.950 5.615 3.610 ;
        RECT 5.405 3.450 5.665 3.610 ;
        RECT 4.445 5.010 4.705 5.170 ;
        RECT 0.175 5.010 4.655 5.170 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.495 5.010 7.055 5.170 ;
        RECT 0.175 5.010 0.815 5.170 ;
  END
END XNR2D1_3
#--------EOF---------

MACRO XOR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.445 4.210 4.705 4.370 ;
        RECT 2.575 4.210 4.655 4.370 ;
        RECT 2.525 4.210 2.785 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 3.450 3.745 3.610 ;
        RECT 3.535 3.450 4.175 3.610 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 2.170 ;
        RECT 2.095 2.010 5.135 2.170 ;
        RECT 4.925 2.010 5.185 2.170 ;
        RECT 2.095 3.450 2.255 5.170 ;
        RECT 2.045 3.450 2.305 3.610 ;
        RECT 2.045 2.010 2.305 2.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 2.575 0.950 3.215 1.110 ;
        RECT 2.575 0.290 2.735 1.110 ;
        RECT 0.655 0.290 2.735 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 3.055 5.010 3.215 5.830 ;
        RECT 0.655 5.670 3.215 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 3.055 0.290 5.135 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 1.615 2.970 2.735 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 2.575 2.970 5.135 3.130 ;
        RECT 4.975 2.970 5.135 5.170 ;
  END
END XOR2D1
MACRO XOR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 3.695 0.450 ;
        RECT 3.485 0.290 3.745 0.450 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 3.215 2.170 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 0.175 0.950 5.135 1.110 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 1.510 ;
        RECT 1.135 1.350 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 1.135 1.350 1.295 5.170 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 2.045 2.490 2.305 2.650 ;
        RECT 2.095 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 5.405 2.490 5.665 2.650 ;
        RECT 5.455 0.290 5.615 2.650 ;
        RECT 4.015 0.290 5.615 0.450 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 1.615 3.450 1.775 5.830 ;
        RECT 0.655 5.670 1.775 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 4.015 2.490 4.175 5.170 ;
  END
END XOR2D1_1
MACRO XOR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 3.695 0.450 ;
        RECT 3.485 0.290 3.745 0.450 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 6.845 5.010 7.105 5.170 ;
        RECT 0.175 0.950 4.655 1.110 ;
        RECT 4.495 0.290 4.655 1.110 ;
        RECT 4.495 0.290 7.055 0.450 ;
        RECT 6.895 0.290 7.055 1.110 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 6.895 0.950 7.055 5.170 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 1.510 ;
        RECT 1.135 1.350 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 1.135 1.350 1.295 5.170 ;
  END
END XOR2D1_2
MACRO XOR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 1.775 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.950 3.695 1.110 ;
        RECT 3.535 0.950 3.695 5.170 ;
        RECT 3.055 5.010 3.695 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 2.095 5.010 2.255 5.830 ;
        RECT 2.095 5.670 6.575 5.830 ;
        RECT 6.365 5.670 6.625 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.085 0.290 1.345 0.450 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 5.010 1.295 5.830 ;
        RECT 1.085 5.670 1.345 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 2.735 2.170 ;
        RECT 2.575 2.010 2.735 3.130 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 4.015 0.950 5.135 1.110 ;
        RECT 4.015 0.950 4.175 3.130 ;
        RECT 3.965 2.970 4.225 3.130 ;
        RECT 4.015 2.970 4.175 4.830 ;
        RECT 4.015 4.670 5.135 4.830 ;
        RECT 4.975 4.670 5.135 5.170 ;
  END
END XOR2D1_3
#--------EOF---------

MACRO XOR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 4.445 4.210 4.705 4.370 ;
        RECT 2.575 4.210 4.655 4.370 ;
        RECT 2.525 4.210 2.785 4.370 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 3.450 3.745 3.610 ;
        RECT 3.535 3.450 4.175 3.610 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.950 2.255 2.170 ;
        RECT 2.095 2.010 5.135 2.170 ;
        RECT 4.925 2.010 5.185 2.170 ;
        RECT 2.095 3.450 2.255 5.170 ;
        RECT 2.045 3.450 2.305 3.610 ;
        RECT 2.045 2.010 2.305 2.170 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 2.575 0.950 3.215 1.110 ;
        RECT 2.575 0.290 2.735 1.110 ;
        RECT 0.655 0.290 2.735 0.450 ;
        RECT 0.605 0.290 0.865 0.450 ;
        RECT 3.055 5.010 3.215 5.830 ;
        RECT 0.655 5.670 3.215 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 3.005 0.290 3.265 0.450 ;
        RECT 3.055 0.290 5.135 0.450 ;
        RECT 4.975 0.290 5.135 1.110 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 1.615 2.970 2.735 3.130 ;
        RECT 1.565 2.970 1.825 3.130 ;
        RECT 2.575 2.970 5.135 3.130 ;
        RECT 4.975 2.970 5.135 5.170 ;
  END
END XOR2D1
MACRO XOR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 3.695 0.450 ;
        RECT 3.485 0.290 3.745 0.450 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 3.215 2.170 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 6.845 4.670 7.105 4.830 ;
        RECT 6.895 0.950 7.055 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 0.175 0.950 5.135 1.110 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 4.975 0.950 5.135 5.170 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 1.510 ;
        RECT 1.135 1.350 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 1.135 1.350 1.295 5.170 ;
        RECT 3.965 0.950 4.225 1.110 ;
        RECT 3.965 5.010 4.225 5.170 ;
        RECT 2.045 2.490 2.305 2.650 ;
        RECT 2.095 2.490 4.655 2.650 ;
        RECT 4.445 2.490 4.705 2.650 ;
        RECT 5.405 2.490 5.665 2.650 ;
        RECT 5.455 0.290 5.615 2.650 ;
        RECT 4.015 0.290 5.615 0.450 ;
        RECT 4.015 0.290 4.175 1.110 ;
        RECT 1.565 3.450 1.825 3.610 ;
        RECT 1.615 3.450 1.775 5.830 ;
        RECT 0.655 5.670 1.775 5.830 ;
        RECT 0.605 5.670 0.865 5.830 ;
        RECT 4.015 2.490 4.175 5.170 ;
  END
END XOR2D1_1
MACRO XOR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.290 2.785 0.450 ;
        RECT 2.575 0.290 3.695 0.450 ;
        RECT 3.485 0.290 3.745 0.450 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.010 2.785 2.170 ;
        RECT 2.575 2.010 2.735 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 4.670 5.185 4.830 ;
        RECT 4.975 0.950 5.135 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.950 0.385 1.110 ;
        RECT 6.845 0.950 7.105 1.110 ;
        RECT 0.125 5.010 0.385 5.170 ;
        RECT 6.845 5.010 7.105 5.170 ;
        RECT 0.175 0.950 4.655 1.110 ;
        RECT 4.495 0.290 4.655 1.110 ;
        RECT 4.495 0.290 7.055 0.450 ;
        RECT 6.895 0.290 7.055 1.110 ;
        RECT 0.175 0.950 0.335 5.170 ;
        RECT 6.895 0.950 7.055 5.170 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.135 0.950 1.295 1.510 ;
        RECT 1.135 1.350 4.655 1.510 ;
        RECT 4.445 1.350 4.705 1.510 ;
        RECT 1.135 1.350 1.295 5.170 ;
  END
END XOR2D1_2
MACRO XOR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.490 1.825 2.650 ;
        RECT 1.615 2.490 1.775 3.130 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.010 0.865 2.170 ;
        RECT 0.655 2.010 0.815 2.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.950 6.145 1.110 ;
        RECT 5.885 4.670 6.145 4.830 ;
        RECT 5.935 0.950 6.095 4.830 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 6.020 7.480 6.220 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.100 7.480 0.100 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.950 3.265 1.110 ;
        RECT 3.005 5.010 3.265 5.170 ;
        RECT 3.055 0.950 3.695 1.110 ;
        RECT 3.535 0.950 3.695 5.170 ;
        RECT 3.055 5.010 3.695 5.170 ;
        RECT 2.045 0.950 2.305 1.110 ;
        RECT 2.045 5.010 2.305 5.170 ;
        RECT 2.095 0.290 2.255 1.110 ;
        RECT 2.095 0.290 6.575 0.450 ;
        RECT 6.365 0.290 6.625 0.450 ;
        RECT 2.095 5.010 2.255 5.830 ;
        RECT 2.095 5.670 6.575 5.830 ;
        RECT 6.365 5.670 6.625 5.830 ;
        RECT 1.085 0.950 1.345 1.110 ;
        RECT 1.085 5.010 1.345 5.170 ;
        RECT 1.085 4.670 1.345 4.830 ;
        RECT 1.135 0.290 1.295 1.110 ;
        RECT 1.085 0.290 1.345 0.450 ;
        RECT 1.135 0.950 1.295 4.830 ;
        RECT 1.135 5.010 1.295 5.830 ;
        RECT 1.085 5.670 1.345 5.830 ;
        RECT 4.925 0.950 5.185 1.110 ;
        RECT 4.925 5.010 5.185 5.170 ;
        RECT 1.565 2.010 1.825 2.170 ;
        RECT 1.615 2.010 2.735 2.170 ;
        RECT 2.575 2.010 2.735 3.130 ;
        RECT 2.525 2.970 2.785 3.130 ;
        RECT 4.015 0.950 5.135 1.110 ;
        RECT 4.015 0.950 4.175 3.130 ;
        RECT 3.965 2.970 4.225 3.130 ;
        RECT 4.015 2.970 4.175 4.830 ;
        RECT 4.015 4.670 5.135 4.830 ;
        RECT 4.975 4.670 5.135 5.170 ;
  END
END XOR2D1_3
#--------EOF---------


END LIBRARY
