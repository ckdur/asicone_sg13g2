VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sg13g2_bpd60
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 60.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 55.930 60.000 60.000 ;
        RECT 0.000 4.070 4.070 55.930 ;
        RECT 55.930 4.070 60.000 55.930 ;
        RECT 0.000 0.000 60.000 4.070 ;
      LAYER Metal4 ;
        RECT 0.000 55.930 60.000 60.000 ;
        RECT 0.000 4.070 4.070 55.930 ;
        RECT 55.930 4.070 60.000 55.930 ;
        RECT 0.000 0.000 60.000 4.070 ;
      LAYER Metal5 ;
        RECT 0.000 55.930 60.000 60.000 ;
        RECT 0.000 4.070 4.070 55.930 ;
        RECT 55.930 4.070 60.000 55.930 ;
        RECT 0.000 0.000 60.000 4.070 ;
      LAYER TopMetal1 ;
        RECT 0.000 55.930 60.000 60.000 ;
        RECT 0.000 4.070 4.070 55.930 ;
        RECT 55.930 4.070 60.000 55.930 ;
        RECT 0.000 0.000 60.000 4.070 ;
      LAYER TopMetal2 ;
        RECT 0.000 57.900 60.000 60.000 ;
        RECT 0.000 57.015 2.985 57.900 ;
        RECT 3.080 57.015 4.980 57.900 ;
        RECT 5.080 57.015 6.980 57.900 ;
        RECT 7.075 57.015 8.975 57.900 ;
        RECT 9.075 57.015 10.975 57.900 ;
        RECT 11.070 57.015 12.970 57.900 ;
        RECT 13.070 57.015 14.970 57.900 ;
        RECT 15.065 57.015 16.965 57.900 ;
        RECT 17.065 57.015 18.965 57.900 ;
        RECT 19.060 57.015 20.960 57.900 ;
        RECT 21.060 57.015 22.960 57.900 ;
        RECT 23.055 57.015 24.955 57.900 ;
        RECT 25.055 57.015 26.955 57.900 ;
        RECT 27.050 57.015 28.950 57.900 ;
        RECT 29.050 57.015 30.950 57.900 ;
        RECT 31.045 57.015 32.945 57.900 ;
        RECT 33.045 57.015 34.945 57.900 ;
        RECT 35.040 57.015 36.940 57.900 ;
        RECT 37.040 57.015 38.940 57.900 ;
        RECT 39.035 57.015 40.935 57.900 ;
        RECT 41.035 57.015 42.935 57.900 ;
        RECT 43.030 57.015 44.930 57.900 ;
        RECT 45.030 57.015 46.930 57.900 ;
        RECT 47.025 57.015 48.925 57.900 ;
        RECT 49.025 57.015 50.925 57.900 ;
        RECT 51.020 57.015 52.920 57.900 ;
        RECT 53.020 57.015 54.920 57.900 ;
        RECT 55.015 57.015 56.915 57.900 ;
        RECT 57.015 57.015 60.000 57.900 ;
        RECT 0.000 56.945 2.100 57.015 ;
        RECT 57.900 56.945 60.000 57.015 ;
        RECT 0.000 55.045 2.985 56.945 ;
        RECT 57.015 55.045 60.000 56.945 ;
        RECT 0.000 54.945 2.100 55.045 ;
        RECT 57.900 54.945 60.000 55.045 ;
        RECT 0.000 53.045 2.985 54.945 ;
        RECT 57.015 53.045 60.000 54.945 ;
        RECT 0.000 52.945 2.100 53.045 ;
        RECT 57.900 52.945 60.000 53.045 ;
        RECT 0.000 51.045 2.985 52.945 ;
        RECT 57.015 51.045 60.000 52.945 ;
        RECT 0.000 50.945 2.100 51.045 ;
        RECT 57.900 50.945 60.000 51.045 ;
        RECT 0.000 49.045 2.985 50.945 ;
        RECT 57.015 49.045 60.000 50.945 ;
        RECT 0.000 48.945 2.100 49.045 ;
        RECT 57.900 48.945 60.000 49.045 ;
        RECT 0.000 47.045 2.985 48.945 ;
        RECT 57.015 47.045 60.000 48.945 ;
        RECT 0.000 46.945 2.100 47.045 ;
        RECT 57.900 46.945 60.000 47.045 ;
        RECT 0.000 45.045 2.985 46.945 ;
        RECT 57.015 45.045 60.000 46.945 ;
        RECT 0.000 44.945 2.100 45.045 ;
        RECT 57.900 44.945 60.000 45.045 ;
        RECT 0.000 43.045 2.985 44.945 ;
        RECT 57.015 43.045 60.000 44.945 ;
        RECT 0.000 42.945 2.100 43.045 ;
        RECT 57.900 42.945 60.000 43.045 ;
        RECT 0.000 41.045 2.985 42.945 ;
        RECT 57.015 41.045 60.000 42.945 ;
        RECT 0.000 40.945 2.100 41.045 ;
        RECT 57.900 40.945 60.000 41.045 ;
        RECT 0.000 39.045 2.985 40.945 ;
        RECT 57.015 39.045 60.000 40.945 ;
        RECT 0.000 38.945 2.100 39.045 ;
        RECT 57.900 38.945 60.000 39.045 ;
        RECT 0.000 37.045 2.985 38.945 ;
        RECT 57.015 37.045 60.000 38.945 ;
        RECT 0.000 36.945 2.100 37.045 ;
        RECT 57.900 36.945 60.000 37.045 ;
        RECT 0.000 35.045 2.985 36.945 ;
        RECT 57.015 35.045 60.000 36.945 ;
        RECT 0.000 34.945 2.100 35.045 ;
        RECT 57.900 34.945 60.000 35.045 ;
        RECT 0.000 33.045 2.985 34.945 ;
        RECT 57.015 33.045 60.000 34.945 ;
        RECT 0.000 32.945 2.100 33.045 ;
        RECT 57.900 32.945 60.000 33.045 ;
        RECT 0.000 31.045 2.985 32.945 ;
        RECT 57.015 31.045 60.000 32.945 ;
        RECT 0.000 30.950 2.100 31.045 ;
        RECT 57.900 30.950 60.000 31.045 ;
        RECT 0.000 29.050 2.985 30.950 ;
        RECT 57.015 29.050 60.000 30.950 ;
        RECT 0.000 28.950 2.100 29.050 ;
        RECT 57.900 28.950 60.000 29.050 ;
        RECT 0.000 27.050 2.985 28.950 ;
        RECT 57.015 27.050 60.000 28.950 ;
        RECT 0.000 26.950 2.100 27.050 ;
        RECT 57.900 26.950 60.000 27.050 ;
        RECT 0.000 25.050 2.985 26.950 ;
        RECT 57.015 25.050 60.000 26.950 ;
        RECT 0.000 24.950 2.100 25.050 ;
        RECT 57.900 24.950 60.000 25.050 ;
        RECT 0.000 23.050 2.985 24.950 ;
        RECT 57.015 23.050 60.000 24.950 ;
        RECT 0.000 22.950 2.100 23.050 ;
        RECT 57.900 22.950 60.000 23.050 ;
        RECT 0.000 21.050 2.985 22.950 ;
        RECT 57.015 21.050 60.000 22.950 ;
        RECT 0.000 20.950 2.100 21.050 ;
        RECT 57.900 20.950 60.000 21.050 ;
        RECT 0.000 19.050 2.985 20.950 ;
        RECT 57.015 19.050 60.000 20.950 ;
        RECT 0.000 18.950 2.100 19.050 ;
        RECT 57.900 18.950 60.000 19.050 ;
        RECT 0.000 17.050 2.985 18.950 ;
        RECT 57.015 17.050 60.000 18.950 ;
        RECT 0.000 16.950 2.100 17.050 ;
        RECT 57.900 16.950 60.000 17.050 ;
        RECT 0.000 15.050 2.985 16.950 ;
        RECT 57.015 15.050 60.000 16.950 ;
        RECT 0.000 14.950 2.100 15.050 ;
        RECT 57.900 14.950 60.000 15.050 ;
        RECT 0.000 13.050 2.985 14.950 ;
        RECT 57.015 13.050 60.000 14.950 ;
        RECT 0.000 12.950 2.100 13.050 ;
        RECT 57.900 12.950 60.000 13.050 ;
        RECT 0.000 11.050 2.985 12.950 ;
        RECT 57.015 11.050 60.000 12.950 ;
        RECT 0.000 10.950 2.100 11.050 ;
        RECT 57.900 10.950 60.000 11.050 ;
        RECT 0.000 9.050 2.985 10.950 ;
        RECT 57.015 9.050 60.000 10.950 ;
        RECT 0.000 8.950 2.100 9.050 ;
        RECT 57.900 8.950 60.000 9.050 ;
        RECT 0.000 7.050 2.985 8.950 ;
        RECT 57.015 7.050 60.000 8.950 ;
        RECT 0.000 6.950 2.100 7.050 ;
        RECT 57.900 6.950 60.000 7.050 ;
        RECT 0.000 5.050 2.985 6.950 ;
        RECT 57.015 5.050 60.000 6.950 ;
        RECT 0.000 4.955 2.100 5.050 ;
        RECT 57.900 4.955 60.000 5.050 ;
        RECT 0.000 3.055 2.985 4.955 ;
        RECT 57.015 3.055 60.000 4.955 ;
        RECT 0.000 2.985 2.100 3.055 ;
        RECT 57.900 2.985 60.000 3.055 ;
        RECT 0.000 2.100 2.985 2.985 ;
        RECT 3.080 2.100 4.980 2.985 ;
        RECT 5.080 2.100 6.980 2.985 ;
        RECT 7.075 2.100 8.975 2.985 ;
        RECT 9.075 2.100 10.975 2.985 ;
        RECT 11.070 2.100 12.970 2.985 ;
        RECT 13.070 2.100 14.970 2.985 ;
        RECT 15.065 2.100 16.965 2.985 ;
        RECT 17.065 2.100 18.965 2.985 ;
        RECT 19.060 2.100 20.960 2.985 ;
        RECT 21.060 2.100 22.960 2.985 ;
        RECT 23.055 2.100 24.955 2.985 ;
        RECT 25.055 2.100 26.955 2.985 ;
        RECT 27.050 2.100 28.950 2.985 ;
        RECT 29.050 2.100 30.950 2.985 ;
        RECT 31.045 2.100 32.945 2.985 ;
        RECT 33.045 2.100 34.945 2.985 ;
        RECT 35.040 2.100 36.940 2.985 ;
        RECT 37.040 2.100 38.940 2.985 ;
        RECT 39.035 2.100 40.935 2.985 ;
        RECT 41.035 2.100 42.935 2.985 ;
        RECT 43.030 2.100 44.930 2.985 ;
        RECT 45.030 2.100 46.930 2.985 ;
        RECT 47.025 2.100 48.925 2.985 ;
        RECT 49.025 2.100 50.925 2.985 ;
        RECT 51.020 2.100 52.920 2.985 ;
        RECT 53.020 2.100 54.920 2.985 ;
        RECT 55.015 2.100 56.915 2.985 ;
        RECT 57.015 2.100 60.000 2.985 ;
        RECT 0.000 0.000 60.000 2.100 ;
  END
END sg13g2_bpd60

#--------EOF---------

MACRO sg13g2_bpd70
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd70 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 70.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 65.930 70.000 70.000 ;
        RECT 0.000 4.070 4.070 65.930 ;
        RECT 65.930 4.070 70.000 65.930 ;
        RECT 0.000 0.000 70.000 4.070 ;
      LAYER Metal4 ;
        RECT 0.000 65.930 70.000 70.000 ;
        RECT 0.000 4.070 4.070 65.930 ;
        RECT 65.930 4.070 70.000 65.930 ;
        RECT 0.000 0.000 70.000 4.070 ;
      LAYER Metal5 ;
        RECT 0.000 65.930 70.000 70.000 ;
        RECT 0.000 4.070 4.070 65.930 ;
        RECT 65.930 4.070 70.000 65.930 ;
        RECT 0.000 0.000 70.000 4.070 ;
      LAYER TopMetal1 ;
        RECT 0.000 65.930 70.000 70.000 ;
        RECT 0.000 4.070 4.070 65.930 ;
        RECT 65.930 4.070 70.000 65.930 ;
        RECT 0.000 0.000 70.000 4.070 ;
      LAYER TopMetal2 ;
        RECT 0.000 67.900 70.000 70.000 ;
        RECT 0.000 67.015 2.985 67.900 ;
        RECT 3.080 67.015 4.980 67.900 ;
        RECT 5.080 67.015 6.980 67.900 ;
        RECT 7.075 67.015 8.975 67.900 ;
        RECT 9.075 67.015 10.975 67.900 ;
        RECT 11.070 67.015 12.970 67.900 ;
        RECT 13.070 67.015 14.970 67.900 ;
        RECT 15.070 67.015 16.970 67.900 ;
        RECT 17.065 67.015 18.965 67.900 ;
        RECT 19.065 67.015 20.965 67.900 ;
        RECT 21.060 67.015 22.960 67.900 ;
        RECT 23.060 67.015 24.960 67.900 ;
        RECT 25.055 67.015 26.955 67.900 ;
        RECT 27.055 67.015 28.955 67.900 ;
        RECT 29.055 67.015 30.955 67.900 ;
        RECT 31.050 67.015 32.950 67.900 ;
        RECT 33.050 67.015 34.950 67.900 ;
        RECT 35.045 67.015 36.945 67.900 ;
        RECT 37.045 67.015 38.945 67.900 ;
        RECT 39.040 67.015 40.940 67.900 ;
        RECT 41.040 67.015 42.940 67.900 ;
        RECT 43.040 67.015 44.940 67.900 ;
        RECT 45.035 67.015 46.935 67.900 ;
        RECT 47.035 67.015 48.935 67.900 ;
        RECT 49.030 67.015 50.930 67.900 ;
        RECT 51.030 67.015 52.930 67.900 ;
        RECT 53.025 67.015 54.925 67.900 ;
        RECT 55.025 67.015 56.925 67.900 ;
        RECT 57.025 67.015 58.925 67.900 ;
        RECT 59.020 67.015 60.920 67.900 ;
        RECT 61.020 67.015 62.920 67.900 ;
        RECT 63.015 67.015 64.915 67.900 ;
        RECT 65.015 67.015 66.915 67.900 ;
        RECT 67.015 67.015 70.000 67.900 ;
        RECT 0.000 66.945 2.100 67.015 ;
        RECT 67.900 66.945 70.000 67.015 ;
        RECT 0.000 65.045 2.985 66.945 ;
        RECT 67.015 65.045 70.000 66.945 ;
        RECT 0.000 64.945 2.100 65.045 ;
        RECT 67.900 64.945 70.000 65.045 ;
        RECT 0.000 63.045 2.985 64.945 ;
        RECT 67.015 63.045 70.000 64.945 ;
        RECT 0.000 62.945 2.100 63.045 ;
        RECT 67.900 62.945 70.000 63.045 ;
        RECT 0.000 61.045 2.985 62.945 ;
        RECT 67.015 61.045 70.000 62.945 ;
        RECT 0.000 60.945 2.100 61.045 ;
        RECT 67.900 60.945 70.000 61.045 ;
        RECT 0.000 59.045 2.985 60.945 ;
        RECT 67.015 59.045 70.000 60.945 ;
        RECT 0.000 58.945 2.100 59.045 ;
        RECT 67.900 58.945 70.000 59.045 ;
        RECT 0.000 57.045 2.985 58.945 ;
        RECT 67.015 57.045 70.000 58.945 ;
        RECT 0.000 56.945 2.100 57.045 ;
        RECT 67.900 56.945 70.000 57.045 ;
        RECT 0.000 55.045 2.985 56.945 ;
        RECT 67.015 55.045 70.000 56.945 ;
        RECT 0.000 54.945 2.100 55.045 ;
        RECT 67.900 54.945 70.000 55.045 ;
        RECT 0.000 53.045 2.985 54.945 ;
        RECT 67.015 53.045 70.000 54.945 ;
        RECT 0.000 52.945 2.100 53.045 ;
        RECT 67.900 52.945 70.000 53.045 ;
        RECT 0.000 51.045 2.985 52.945 ;
        RECT 67.015 51.045 70.000 52.945 ;
        RECT 0.000 50.945 2.100 51.045 ;
        RECT 67.900 50.945 70.000 51.045 ;
        RECT 0.000 49.045 2.985 50.945 ;
        RECT 67.015 49.045 70.000 50.945 ;
        RECT 0.000 48.945 2.100 49.045 ;
        RECT 67.900 48.945 70.000 49.045 ;
        RECT 0.000 47.045 2.985 48.945 ;
        RECT 67.015 47.045 70.000 48.945 ;
        RECT 0.000 46.945 2.100 47.045 ;
        RECT 67.900 46.945 70.000 47.045 ;
        RECT 0.000 45.045 2.985 46.945 ;
        RECT 67.015 45.045 70.000 46.945 ;
        RECT 0.000 44.945 2.100 45.045 ;
        RECT 67.900 44.945 70.000 45.045 ;
        RECT 0.000 43.045 2.985 44.945 ;
        RECT 67.015 43.045 70.000 44.945 ;
        RECT 0.000 42.945 2.100 43.045 ;
        RECT 67.900 42.945 70.000 43.045 ;
        RECT 0.000 41.045 2.985 42.945 ;
        RECT 67.015 41.045 70.000 42.945 ;
        RECT 0.000 40.945 2.100 41.045 ;
        RECT 67.900 40.945 70.000 41.045 ;
        RECT 0.000 39.045 2.985 40.945 ;
        RECT 67.015 39.045 70.000 40.945 ;
        RECT 0.000 38.945 2.100 39.045 ;
        RECT 67.900 38.945 70.000 39.045 ;
        RECT 0.000 37.045 2.985 38.945 ;
        RECT 67.015 37.045 70.000 38.945 ;
        RECT 0.000 36.945 2.100 37.045 ;
        RECT 67.900 36.945 70.000 37.045 ;
        RECT 0.000 35.045 2.985 36.945 ;
        RECT 67.015 35.045 70.000 36.945 ;
        RECT 0.000 34.950 2.100 35.045 ;
        RECT 67.900 34.950 70.000 35.045 ;
        RECT 0.000 33.050 2.985 34.950 ;
        RECT 67.015 33.050 70.000 34.950 ;
        RECT 0.000 32.950 2.100 33.050 ;
        RECT 67.900 32.950 70.000 33.050 ;
        RECT 0.000 31.050 2.985 32.950 ;
        RECT 67.015 31.050 70.000 32.950 ;
        RECT 0.000 30.950 2.100 31.050 ;
        RECT 67.900 30.950 70.000 31.050 ;
        RECT 0.000 29.050 2.985 30.950 ;
        RECT 67.015 29.050 70.000 30.950 ;
        RECT 0.000 28.950 2.100 29.050 ;
        RECT 67.900 28.950 70.000 29.050 ;
        RECT 0.000 27.050 2.985 28.950 ;
        RECT 67.015 27.050 70.000 28.950 ;
        RECT 0.000 26.950 2.100 27.050 ;
        RECT 67.900 26.950 70.000 27.050 ;
        RECT 0.000 25.050 2.985 26.950 ;
        RECT 67.015 25.050 70.000 26.950 ;
        RECT 0.000 24.950 2.100 25.050 ;
        RECT 67.900 24.950 70.000 25.050 ;
        RECT 0.000 23.050 2.985 24.950 ;
        RECT 67.015 23.050 70.000 24.950 ;
        RECT 0.000 22.950 2.100 23.050 ;
        RECT 67.900 22.950 70.000 23.050 ;
        RECT 0.000 21.050 2.985 22.950 ;
        RECT 67.015 21.050 70.000 22.950 ;
        RECT 0.000 20.950 2.100 21.050 ;
        RECT 67.900 20.950 70.000 21.050 ;
        RECT 0.000 19.050 2.985 20.950 ;
        RECT 67.015 19.050 70.000 20.950 ;
        RECT 0.000 18.950 2.100 19.050 ;
        RECT 67.900 18.950 70.000 19.050 ;
        RECT 0.000 17.050 2.985 18.950 ;
        RECT 67.015 17.050 70.000 18.950 ;
        RECT 0.000 16.950 2.100 17.050 ;
        RECT 67.900 16.950 70.000 17.050 ;
        RECT 0.000 15.050 2.985 16.950 ;
        RECT 67.015 15.050 70.000 16.950 ;
        RECT 0.000 14.950 2.100 15.050 ;
        RECT 67.900 14.950 70.000 15.050 ;
        RECT 0.000 13.050 2.985 14.950 ;
        RECT 67.015 13.050 70.000 14.950 ;
        RECT 0.000 12.950 2.100 13.050 ;
        RECT 67.900 12.950 70.000 13.050 ;
        RECT 0.000 11.050 2.985 12.950 ;
        RECT 67.015 11.050 70.000 12.950 ;
        RECT 0.000 10.950 2.100 11.050 ;
        RECT 67.900 10.950 70.000 11.050 ;
        RECT 0.000 9.050 2.985 10.950 ;
        RECT 67.015 9.050 70.000 10.950 ;
        RECT 0.000 8.950 2.100 9.050 ;
        RECT 67.900 8.950 70.000 9.050 ;
        RECT 0.000 7.050 2.985 8.950 ;
        RECT 67.015 7.050 70.000 8.950 ;
        RECT 0.000 6.950 2.100 7.050 ;
        RECT 67.900 6.950 70.000 7.050 ;
        RECT 0.000 5.050 2.985 6.950 ;
        RECT 67.015 5.050 70.000 6.950 ;
        RECT 0.000 4.955 2.100 5.050 ;
        RECT 67.900 4.955 70.000 5.050 ;
        RECT 0.000 3.055 2.985 4.955 ;
        RECT 67.015 3.055 70.000 4.955 ;
        RECT 0.000 2.985 2.100 3.055 ;
        RECT 67.900 2.985 70.000 3.055 ;
        RECT 0.000 2.100 2.985 2.985 ;
        RECT 3.080 2.100 4.980 2.985 ;
        RECT 5.080 2.100 6.980 2.985 ;
        RECT 7.075 2.100 8.975 2.985 ;
        RECT 9.075 2.100 10.975 2.985 ;
        RECT 11.070 2.100 12.970 2.985 ;
        RECT 13.070 2.100 14.970 2.985 ;
        RECT 15.070 2.100 16.970 2.985 ;
        RECT 17.065 2.100 18.965 2.985 ;
        RECT 19.065 2.100 20.965 2.985 ;
        RECT 21.060 2.100 22.960 2.985 ;
        RECT 23.060 2.100 24.960 2.985 ;
        RECT 25.055 2.100 26.955 2.985 ;
        RECT 27.055 2.100 28.955 2.985 ;
        RECT 29.055 2.100 30.955 2.985 ;
        RECT 31.050 2.100 32.950 2.985 ;
        RECT 33.050 2.100 34.950 2.985 ;
        RECT 35.045 2.100 36.945 2.985 ;
        RECT 37.045 2.100 38.945 2.985 ;
        RECT 39.040 2.100 40.940 2.985 ;
        RECT 41.040 2.100 42.940 2.985 ;
        RECT 43.040 2.100 44.940 2.985 ;
        RECT 45.035 2.100 46.935 2.985 ;
        RECT 47.035 2.100 48.935 2.985 ;
        RECT 49.030 2.100 50.930 2.985 ;
        RECT 51.030 2.100 52.930 2.985 ;
        RECT 53.025 2.100 54.925 2.985 ;
        RECT 55.025 2.100 56.925 2.985 ;
        RECT 57.025 2.100 58.925 2.985 ;
        RECT 59.020 2.100 60.920 2.985 ;
        RECT 61.020 2.100 62.920 2.985 ;
        RECT 63.015 2.100 64.915 2.985 ;
        RECT 65.015 2.100 66.915 2.985 ;
        RECT 67.015 2.100 70.000 2.985 ;
        RECT 0.000 0.000 70.000 2.100 ;
  END
END sg13g2_bpd70

#--------EOF---------

MACRO sg13g2_bpd80
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd80 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 80.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 75.930 80.000 80.000 ;
        RECT 0.000 4.070 4.070 75.930 ;
        RECT 75.930 4.070 80.000 75.930 ;
        RECT 0.000 0.000 80.000 4.070 ;
      LAYER Metal4 ;
        RECT 0.000 75.930 80.000 80.000 ;
        RECT 0.000 4.070 4.070 75.930 ;
        RECT 75.930 4.070 80.000 75.930 ;
        RECT 0.000 0.000 80.000 4.070 ;
      LAYER Metal5 ;
        RECT 0.000 75.930 80.000 80.000 ;
        RECT 0.000 4.070 4.070 75.930 ;
        RECT 75.930 4.070 80.000 75.930 ;
        RECT 0.000 0.000 80.000 4.070 ;
      LAYER TopMetal1 ;
        RECT 0.000 75.930 80.000 80.000 ;
        RECT 0.000 4.070 4.070 75.930 ;
        RECT 75.930 4.070 80.000 75.930 ;
        RECT 0.000 0.000 80.000 4.070 ;
      LAYER TopMetal2 ;
        RECT 0.000 77.900 80.000 80.000 ;
        RECT 0.000 77.015 2.985 77.900 ;
        RECT 3.080 77.015 4.980 77.900 ;
        RECT 5.080 77.015 6.980 77.900 ;
        RECT 7.075 77.015 8.975 77.900 ;
        RECT 9.075 77.015 10.975 77.900 ;
        RECT 11.075 77.015 12.975 77.900 ;
        RECT 13.070 77.015 14.970 77.900 ;
        RECT 15.070 77.015 16.970 77.900 ;
        RECT 17.070 77.015 18.970 77.900 ;
        RECT 19.065 77.015 20.965 77.900 ;
        RECT 21.065 77.015 22.965 77.900 ;
        RECT 23.060 77.015 24.960 77.900 ;
        RECT 25.060 77.015 26.960 77.900 ;
        RECT 27.060 77.015 28.960 77.900 ;
        RECT 29.055 77.015 30.955 77.900 ;
        RECT 31.055 77.015 32.955 77.900 ;
        RECT 33.055 77.015 34.955 77.900 ;
        RECT 35.050 77.015 36.950 77.900 ;
        RECT 37.050 77.015 38.950 77.900 ;
        RECT 39.050 77.015 40.950 77.900 ;
        RECT 41.045 77.015 42.945 77.900 ;
        RECT 43.045 77.015 44.945 77.900 ;
        RECT 45.040 77.015 46.940 77.900 ;
        RECT 47.040 77.015 48.940 77.900 ;
        RECT 49.040 77.015 50.940 77.900 ;
        RECT 51.035 77.015 52.935 77.900 ;
        RECT 53.035 77.015 54.935 77.900 ;
        RECT 55.035 77.015 56.935 77.900 ;
        RECT 57.030 77.015 58.930 77.900 ;
        RECT 59.030 77.015 60.930 77.900 ;
        RECT 61.025 77.015 62.925 77.900 ;
        RECT 63.025 77.015 64.925 77.900 ;
        RECT 65.025 77.015 66.925 77.900 ;
        RECT 67.020 77.015 68.920 77.900 ;
        RECT 69.020 77.015 70.920 77.900 ;
        RECT 71.020 77.015 72.920 77.900 ;
        RECT 73.015 77.015 74.915 77.900 ;
        RECT 75.015 77.015 76.915 77.900 ;
        RECT 77.015 77.015 80.000 77.900 ;
        RECT 0.000 76.945 2.100 77.015 ;
        RECT 77.900 76.945 80.000 77.015 ;
        RECT 0.000 75.045 2.985 76.945 ;
        RECT 77.015 75.045 80.000 76.945 ;
        RECT 0.000 74.945 2.100 75.045 ;
        RECT 77.900 74.945 80.000 75.045 ;
        RECT 0.000 73.045 2.985 74.945 ;
        RECT 77.015 73.045 80.000 74.945 ;
        RECT 0.000 72.945 2.100 73.045 ;
        RECT 77.900 72.945 80.000 73.045 ;
        RECT 0.000 71.045 2.985 72.945 ;
        RECT 77.015 71.045 80.000 72.945 ;
        RECT 0.000 70.945 2.100 71.045 ;
        RECT 77.900 70.945 80.000 71.045 ;
        RECT 0.000 69.045 2.985 70.945 ;
        RECT 77.015 69.045 80.000 70.945 ;
        RECT 0.000 68.945 2.100 69.045 ;
        RECT 77.900 68.945 80.000 69.045 ;
        RECT 0.000 67.045 2.985 68.945 ;
        RECT 77.015 67.045 80.000 68.945 ;
        RECT 0.000 66.945 2.100 67.045 ;
        RECT 77.900 66.945 80.000 67.045 ;
        RECT 0.000 65.045 2.985 66.945 ;
        RECT 77.015 65.045 80.000 66.945 ;
        RECT 0.000 64.945 2.100 65.045 ;
        RECT 77.900 64.945 80.000 65.045 ;
        RECT 0.000 63.045 2.985 64.945 ;
        RECT 77.015 63.045 80.000 64.945 ;
        RECT 0.000 62.945 2.100 63.045 ;
        RECT 77.900 62.945 80.000 63.045 ;
        RECT 0.000 61.045 2.985 62.945 ;
        RECT 77.015 61.045 80.000 62.945 ;
        RECT 0.000 60.945 2.100 61.045 ;
        RECT 77.900 60.945 80.000 61.045 ;
        RECT 0.000 59.045 2.985 60.945 ;
        RECT 77.015 59.045 80.000 60.945 ;
        RECT 0.000 58.945 2.100 59.045 ;
        RECT 77.900 58.945 80.000 59.045 ;
        RECT 0.000 57.045 2.985 58.945 ;
        RECT 77.015 57.045 80.000 58.945 ;
        RECT 0.000 56.945 2.100 57.045 ;
        RECT 77.900 56.945 80.000 57.045 ;
        RECT 0.000 55.045 2.985 56.945 ;
        RECT 77.015 55.045 80.000 56.945 ;
        RECT 0.000 54.945 2.100 55.045 ;
        RECT 77.900 54.945 80.000 55.045 ;
        RECT 0.000 53.045 2.985 54.945 ;
        RECT 77.015 53.045 80.000 54.945 ;
        RECT 0.000 52.945 2.100 53.045 ;
        RECT 77.900 52.945 80.000 53.045 ;
        RECT 0.000 51.045 2.985 52.945 ;
        RECT 77.015 51.045 80.000 52.945 ;
        RECT 0.000 50.945 2.100 51.045 ;
        RECT 77.900 50.945 80.000 51.045 ;
        RECT 0.000 49.045 2.985 50.945 ;
        RECT 77.015 49.045 80.000 50.945 ;
        RECT 0.000 48.945 2.100 49.045 ;
        RECT 77.900 48.945 80.000 49.045 ;
        RECT 0.000 47.045 2.985 48.945 ;
        RECT 77.015 47.045 80.000 48.945 ;
        RECT 0.000 46.945 2.100 47.045 ;
        RECT 77.900 46.945 80.000 47.045 ;
        RECT 0.000 45.045 2.985 46.945 ;
        RECT 77.015 45.045 80.000 46.945 ;
        RECT 0.000 44.945 2.100 45.045 ;
        RECT 77.900 44.945 80.000 45.045 ;
        RECT 0.000 43.045 2.985 44.945 ;
        RECT 77.015 43.045 80.000 44.945 ;
        RECT 0.000 42.945 2.100 43.045 ;
        RECT 77.900 42.945 80.000 43.045 ;
        RECT 0.000 41.045 2.985 42.945 ;
        RECT 77.015 41.045 80.000 42.945 ;
        RECT 0.000 40.950 2.100 41.045 ;
        RECT 77.900 40.950 80.000 41.045 ;
        RECT 0.000 39.050 2.985 40.950 ;
        RECT 77.015 39.050 80.000 40.950 ;
        RECT 0.000 38.950 2.100 39.050 ;
        RECT 77.900 38.950 80.000 39.050 ;
        RECT 0.000 37.050 2.985 38.950 ;
        RECT 77.015 37.050 80.000 38.950 ;
        RECT 0.000 36.950 2.100 37.050 ;
        RECT 77.900 36.950 80.000 37.050 ;
        RECT 0.000 35.050 2.985 36.950 ;
        RECT 77.015 35.050 80.000 36.950 ;
        RECT 0.000 34.950 2.100 35.050 ;
        RECT 77.900 34.950 80.000 35.050 ;
        RECT 0.000 33.050 2.985 34.950 ;
        RECT 77.015 33.050 80.000 34.950 ;
        RECT 0.000 32.950 2.100 33.050 ;
        RECT 77.900 32.950 80.000 33.050 ;
        RECT 0.000 31.050 2.985 32.950 ;
        RECT 77.015 31.050 80.000 32.950 ;
        RECT 0.000 30.950 2.100 31.050 ;
        RECT 77.900 30.950 80.000 31.050 ;
        RECT 0.000 29.050 2.985 30.950 ;
        RECT 77.015 29.050 80.000 30.950 ;
        RECT 0.000 28.950 2.100 29.050 ;
        RECT 77.900 28.950 80.000 29.050 ;
        RECT 0.000 27.050 2.985 28.950 ;
        RECT 77.015 27.050 80.000 28.950 ;
        RECT 0.000 26.950 2.100 27.050 ;
        RECT 77.900 26.950 80.000 27.050 ;
        RECT 0.000 25.050 2.985 26.950 ;
        RECT 77.015 25.050 80.000 26.950 ;
        RECT 0.000 24.950 2.100 25.050 ;
        RECT 77.900 24.950 80.000 25.050 ;
        RECT 0.000 23.050 2.985 24.950 ;
        RECT 77.015 23.050 80.000 24.950 ;
        RECT 0.000 22.950 2.100 23.050 ;
        RECT 77.900 22.950 80.000 23.050 ;
        RECT 0.000 21.050 2.985 22.950 ;
        RECT 77.015 21.050 80.000 22.950 ;
        RECT 0.000 20.950 2.100 21.050 ;
        RECT 77.900 20.950 80.000 21.050 ;
        RECT 0.000 19.050 2.985 20.950 ;
        RECT 77.015 19.050 80.000 20.950 ;
        RECT 0.000 18.950 2.100 19.050 ;
        RECT 77.900 18.950 80.000 19.050 ;
        RECT 0.000 17.050 2.985 18.950 ;
        RECT 77.015 17.050 80.000 18.950 ;
        RECT 0.000 16.950 2.100 17.050 ;
        RECT 77.900 16.950 80.000 17.050 ;
        RECT 0.000 15.050 2.985 16.950 ;
        RECT 77.015 15.050 80.000 16.950 ;
        RECT 0.000 14.950 2.100 15.050 ;
        RECT 77.900 14.950 80.000 15.050 ;
        RECT 0.000 13.050 2.985 14.950 ;
        RECT 77.015 13.050 80.000 14.950 ;
        RECT 0.000 12.950 2.100 13.050 ;
        RECT 77.900 12.950 80.000 13.050 ;
        RECT 0.000 11.050 2.985 12.950 ;
        RECT 77.015 11.050 80.000 12.950 ;
        RECT 0.000 10.950 2.100 11.050 ;
        RECT 77.900 10.950 80.000 11.050 ;
        RECT 0.000 9.050 2.985 10.950 ;
        RECT 77.015 9.050 80.000 10.950 ;
        RECT 0.000 8.950 2.100 9.050 ;
        RECT 77.900 8.950 80.000 9.050 ;
        RECT 0.000 7.050 2.985 8.950 ;
        RECT 77.015 7.050 80.000 8.950 ;
        RECT 0.000 6.950 2.100 7.050 ;
        RECT 77.900 6.950 80.000 7.050 ;
        RECT 0.000 5.050 2.985 6.950 ;
        RECT 77.015 5.050 80.000 6.950 ;
        RECT 0.000 4.955 2.100 5.050 ;
        RECT 77.900 4.955 80.000 5.050 ;
        RECT 0.000 3.055 2.985 4.955 ;
        RECT 77.015 3.055 80.000 4.955 ;
        RECT 0.000 2.985 2.100 3.055 ;
        RECT 77.900 2.985 80.000 3.055 ;
        RECT 0.000 2.100 2.985 2.985 ;
        RECT 3.080 2.100 4.980 2.985 ;
        RECT 5.080 2.100 6.980 2.985 ;
        RECT 7.075 2.100 8.975 2.985 ;
        RECT 9.075 2.100 10.975 2.985 ;
        RECT 11.075 2.100 12.975 2.985 ;
        RECT 13.070 2.100 14.970 2.985 ;
        RECT 15.070 2.100 16.970 2.985 ;
        RECT 17.070 2.100 18.970 2.985 ;
        RECT 19.065 2.100 20.965 2.985 ;
        RECT 21.065 2.100 22.965 2.985 ;
        RECT 23.060 2.100 24.960 2.985 ;
        RECT 25.060 2.100 26.960 2.985 ;
        RECT 27.060 2.100 28.960 2.985 ;
        RECT 29.055 2.100 30.955 2.985 ;
        RECT 31.055 2.100 32.955 2.985 ;
        RECT 33.055 2.100 34.955 2.985 ;
        RECT 35.050 2.100 36.950 2.985 ;
        RECT 37.050 2.100 38.950 2.985 ;
        RECT 39.050 2.100 40.950 2.985 ;
        RECT 41.045 2.100 42.945 2.985 ;
        RECT 43.045 2.100 44.945 2.985 ;
        RECT 45.040 2.100 46.940 2.985 ;
        RECT 47.040 2.100 48.940 2.985 ;
        RECT 49.040 2.100 50.940 2.985 ;
        RECT 51.035 2.100 52.935 2.985 ;
        RECT 53.035 2.100 54.935 2.985 ;
        RECT 55.035 2.100 56.935 2.985 ;
        RECT 57.030 2.100 58.930 2.985 ;
        RECT 59.030 2.100 60.930 2.985 ;
        RECT 61.025 2.100 62.925 2.985 ;
        RECT 63.025 2.100 64.925 2.985 ;
        RECT 65.025 2.100 66.925 2.985 ;
        RECT 67.020 2.100 68.920 2.985 ;
        RECT 69.020 2.100 70.920 2.985 ;
        RECT 71.020 2.100 72.920 2.985 ;
        RECT 73.015 2.100 74.915 2.985 ;
        RECT 75.015 2.100 76.915 2.985 ;
        RECT 77.015 2.100 80.000 2.985 ;
        RECT 0.000 0.000 80.000 2.100 ;
  END
END sg13g2_bpd80

#--------EOF---------


END LIBRARY
