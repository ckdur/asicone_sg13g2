VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.34 BY 6.12 ;
END obssite

#--------EOF---------

MACRO AN2D0
  CLASS CORE ;
  FOREIGN AN2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN z
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 1.150 3.215 4.970 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a2
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 1.630 2.215 1.760 4.600 ;
        RECT 1.065 2.085 1.760 2.215 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 1.630 1.280 1.760 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.135 2.230 1.295 2.710 ;
        RECT 1.085 2.070 1.345 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.970 1.775 5.130 ;
        RECT 1.615 2.230 1.775 4.970 ;
        RECT 1.615 2.070 2.785 2.230 ;
        RECT 1.615 1.150 1.775 2.070 ;
        RECT 0.125 0.990 1.775 1.150 ;
  END
END AN2D0

#--------EOF---------

MACRO AN2D1
  CLASS CORE ;
  FOREIGN AN2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.241150 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.575 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 3.005 1.410 3.265 1.570 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.241150 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 1.065 2.085 1.760 2.215 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 1.630 1.575 1.760 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.135 2.230 1.295 2.710 ;
        RECT 1.085 2.070 1.345 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 1.775 4.230 ;
        RECT 1.615 2.230 1.775 4.070 ;
        RECT 1.615 2.070 2.785 2.230 ;
        RECT 1.615 1.150 1.775 2.070 ;
        RECT 0.125 0.990 1.775 1.150 ;
  END
END AN2D1

#--------EOF---------

MACRO AN2D2
  CLASS CORE ;
  FOREIGN AN2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 0.670 2.085 1.845 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 1.615 1.570 1.775 2.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.615 1.410 4.225 1.570 ;
  END
END AN2D2

#--------EOF---------

MACRO AN2D4
  CLASS CORE ;
  FOREIGN AN2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 2.780 1.760 4.000 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 2.215 1.760 2.480 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 1.630 2.085 2.720 2.215 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.550 2.255 2.710 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 4.925 1.410 7.105 1.570 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 2.985 2.215 3.285 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 2.985 2.085 3.680 2.215 ;
        RECT 2.985 2.000 3.285 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 0.605 2.070 3.265 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 3.945 3.175 4.245 3.260 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 3.945 3.045 4.640 3.175 ;
        RECT 3.945 2.960 4.245 3.045 ;
        RECT 4.510 2.300 4.640 3.045 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 4.425 2.085 7.520 2.215 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.135 3.190 1.295 4.070 ;
        RECT 3.055 3.190 3.215 4.070 ;
        RECT 1.135 3.030 4.225 3.190 ;
        RECT 4.445 2.070 4.705 2.230 ;
        RECT 4.495 1.570 4.655 2.070 ;
        RECT 2.045 1.410 4.655 1.570 ;
  END
END AN2D4

#--------EOF---------

MACRO AO21D0
  CLASS CORE ;
  FOREIGN AO21D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.600 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.280 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.780 1.760 4.600 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 1.280 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.710 1.775 3.190 ;
        RECT 1.565 2.550 1.825 2.710 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 5.630 3.695 5.790 ;
        RECT 2.575 5.130 2.735 5.630 ;
        RECT 3.535 5.130 3.695 5.630 ;
        RECT 2.045 4.970 2.735 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 2.095 2.230 2.255 4.630 ;
        RECT 0.605 2.070 2.255 2.230 ;
        RECT 2.095 1.150 2.255 2.070 ;
        RECT 2.045 0.990 2.305 1.150 ;
  END
END AO21D0

#--------EOF---------

MACRO AO21D1
  CLASS CORE ;
  FOREIGN AO21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.780 1.760 4.000 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 1.640 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.710 1.775 3.190 ;
        RECT 1.565 2.550 1.825 2.710 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 4.225 4.790 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 3.055 3.190 3.215 4.070 ;
        RECT 2.095 3.030 3.215 3.190 ;
        RECT 2.095 2.230 2.255 3.030 ;
        RECT 0.605 2.070 2.255 2.230 ;
        RECT 2.095 1.570 2.255 2.070 ;
        RECT 2.045 1.410 2.305 1.570 ;
  END
END AO21D1

#--------EOF---------

MACRO AO21D2
  CLASS CORE ;
  FOREIGN AO21D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.000 4.725 2.300 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.780 2.720 4.000 ;
        RECT 2.505 2.480 2.805 2.780 ;
        RECT 2.590 1.640 2.720 2.480 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.710 2.735 3.190 ;
        RECT 2.525 2.550 2.785 2.710 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 0.670 2.085 1.845 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 4.630 5.185 4.790 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 4.015 3.190 4.175 4.070 ;
        RECT 3.055 3.030 4.175 3.190 ;
        RECT 3.055 2.230 3.215 3.030 ;
        RECT 1.565 2.070 3.215 2.230 ;
        RECT 3.055 1.570 3.215 2.070 ;
        RECT 3.005 1.410 3.265 1.570 ;
  END
END AO21D2

#--------EOF---------

MACRO AO21D4
  CLASS CORE ;
  FOREIGN AO21D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.540 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 0.585 2.085 5.600 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 3.260 1.760 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 1.545 2.960 1.845 3.260 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 1.545 0.475 1.845 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 1.545 0.345 4.640 0.475 ;
        RECT 1.545 0.260 1.845 0.345 ;
      LAYER Metal1 ;
        RECT 1.565 3.030 4.705 3.190 ;
        RECT 1.615 0.490 1.775 3.030 ;
        RECT 1.565 0.330 1.825 0.490 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
      LAYER Metal1 ;
        RECT 0.655 3.190 0.815 4.230 ;
        RECT 0.605 3.030 0.865 3.190 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 8.815 1.570 8.975 4.070 ;
        RECT 6.845 1.410 9.025 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 0.000 -0.150 10.540 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 10.540 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 5.470 3.820 5.600 4.000 ;
        RECT 6.430 2.300 6.560 4.000 ;
        RECT 6.345 2.215 6.645 2.300 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 6.345 2.085 9.440 2.215 ;
        RECT 6.345 2.000 6.645 2.085 ;
        RECT 2.590 1.640 2.720 1.820 ;
        RECT 3.550 1.640 3.680 1.820 ;
        RECT 6.430 1.640 6.560 2.000 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.630 5.185 4.790 ;
        RECT 2.045 4.070 5.135 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 6.365 2.070 6.625 2.230 ;
        RECT 6.415 1.570 6.575 2.070 ;
        RECT 2.045 1.410 6.575 1.570 ;
  END
END AO21D4

#--------EOF---------

MACRO AOI21D0
  CLASS CORE ;
  FOREIGN AOI21D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.796800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 1.135 4.630 2.255 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.655 5.630 1.775 5.790 ;
        RECT 0.655 5.130 0.815 5.630 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 1.615 5.130 1.775 5.630 ;
        RECT 1.615 4.970 2.305 5.130 ;
  END
END AOI21D0

#--------EOF---------

MACRO AOI21D1
  CLASS CORE ;
  FOREIGN AOI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 3.190 1.295 4.070 ;
        RECT 1.135 3.030 2.255 3.190 ;
        RECT 2.095 1.570 2.255 3.030 ;
        RECT 2.045 1.410 2.305 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 2.305 4.790 ;
  END
END AOI21D1

#--------EOF---------

MACRO AOI21D2
  CLASS CORE ;
  FOREIGN AOI21D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 2.045 1.410 4.225 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 1.545 2.085 4.640 2.215 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 3.260 2.720 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 2.505 2.960 2.805 3.260 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 0.670 1.640 0.800 2.960 ;
        RECT 5.470 1.640 5.600 3.045 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 0.670 0.345 5.600 0.475 ;
      LAYER Metal1 ;
        RECT 0.655 4.630 2.735 4.790 ;
        RECT 0.655 3.190 0.815 4.630 ;
        RECT 2.575 3.190 2.735 4.630 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 2.525 3.030 2.785 3.190 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.585 5.560 0.885 5.860 ;
        RECT 0.670 5.200 0.800 5.560 ;
        RECT 0.670 3.820 0.800 4.000 ;
      LAYER Metal1 ;
        RECT 0.605 5.630 0.865 5.790 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 5.470 3.820 5.600 4.000 ;
        RECT 2.590 1.640 2.720 1.820 ;
        RECT 3.550 1.640 3.680 1.820 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.970 3.215 5.130 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 3.005 4.630 5.185 4.790 ;
  END
END AOI21D2

#--------EOF---------

MACRO AOI21D4
  CLASS CORE ;
  FOREIGN AOI21D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.374400 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 10.685 4.070 10.945 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 8.815 1.570 8.975 4.070 ;
        RECT 10.735 1.570 10.895 4.070 ;
        RECT 4.925 1.410 10.945 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 5.385 2.215 5.685 2.300 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 4.510 2.085 11.360 2.215 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.385 2.000 5.685 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
      LAYER Metal1 ;
        RECT 5.455 2.230 5.615 2.710 ;
        RECT 5.405 2.070 5.665 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 2.590 3.260 2.720 4.000 ;
        RECT 2.505 3.175 2.805 3.260 ;
        RECT 3.550 3.175 3.680 4.000 ;
        RECT 0.670 3.045 3.680 3.175 ;
        RECT 2.505 2.960 2.805 3.045 ;
        RECT 5.470 1.640 5.600 1.820 ;
        RECT 6.430 1.640 6.560 1.820 ;
        RECT 9.310 1.640 9.440 1.820 ;
        RECT 10.270 1.640 10.400 1.820 ;
        RECT 4.425 0.475 4.725 0.560 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 6.430 0.475 6.560 0.920 ;
        RECT 9.310 0.475 9.440 0.920 ;
        RECT 10.270 0.475 10.400 0.920 ;
        RECT 4.425 0.345 10.400 0.475 ;
        RECT 4.425 0.260 4.725 0.345 ;
      LAYER Metal1 ;
        RECT 2.525 3.030 2.785 3.190 ;
        RECT 2.575 2.230 2.735 3.030 ;
        RECT 2.575 2.070 4.655 2.230 ;
        RECT 4.495 0.490 4.655 2.070 ;
        RECT 4.445 0.330 4.705 0.490 ;
    END
  END b
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 4.510 2.695 4.640 4.000 ;
        RECT 5.470 2.695 5.600 4.000 ;
        RECT 7.390 3.175 7.520 4.000 ;
        RECT 8.350 3.260 8.480 4.000 ;
        RECT 8.265 3.175 8.565 3.260 ;
        RECT 7.390 3.045 8.565 3.175 ;
        RECT 8.265 2.960 8.565 3.045 ;
        RECT 5.865 2.695 6.165 2.780 ;
        RECT 4.030 2.565 6.165 2.695 ;
        RECT 4.030 2.215 4.160 2.565 ;
        RECT 5.865 2.480 6.165 2.565 ;
        RECT 0.670 2.085 4.160 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 6.415 4.630 8.495 4.790 ;
        RECT 6.415 2.710 6.575 4.630 ;
        RECT 8.335 3.190 8.495 4.630 ;
        RECT 8.285 3.030 8.545 3.190 ;
        RECT 5.885 2.550 6.575 2.710 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 4.015 5.630 11.855 5.790 ;
        RECT 4.015 5.130 4.175 5.630 ;
        RECT 5.935 5.130 6.095 5.630 ;
        RECT 7.855 5.130 8.015 5.630 ;
        RECT 9.775 5.130 9.935 5.630 ;
        RECT 11.695 5.130 11.855 5.630 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 4.495 4.970 11.375 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
        RECT 3.535 4.790 3.695 4.970 ;
        RECT 0.125 4.630 3.695 4.790 ;
        RECT 4.495 4.230 4.655 4.970 ;
        RECT 2.095 4.070 4.655 4.230 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 11.215 1.570 11.375 4.970 ;
        RECT 0.125 1.410 3.695 1.570 ;
        RECT 11.215 1.410 11.905 1.570 ;
        RECT 2.095 1.150 2.255 1.410 ;
        RECT 3.535 1.150 3.695 1.410 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.535 0.990 4.225 1.150 ;
  END
END AOI21D4

#--------EOF---------

MACRO ANTENNA
  CLASS CORE ANTENNACELL ;
  FOREIGN ANTENNA ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.380 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.380 6.270 ;
    END
  END vdd
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.440450 ;
    ANTENNADIFFAREA 2.880900 ;
    PORT
      LAYER Metal1 ;
        RECT 0.590 5.040 1.810 5.200 ;
        RECT 0.640 1.080 0.800 5.040 ;
        RECT 0.590 0.920 1.810 1.080 ;
    END
  END i
END ANTENNA

#--------EOF---------

MACRO BUFFD0
  CLASS CORE ;
  FOREIGN BUFFD0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.486775 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 1.150 2.255 4.970 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.078650 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.840 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.165 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.065 1.555 1.365 1.640 ;
        RECT 1.630 1.555 1.760 4.615 ;
        RECT 1.065 1.425 1.760 1.555 ;
        RECT 1.065 1.340 1.365 1.425 ;
        RECT 1.630 1.170 1.760 1.425 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 1.570 0.335 4.970 ;
        RECT 0.175 1.410 1.345 1.570 ;
        RECT 0.175 1.150 0.335 1.410 ;
        RECT 0.125 0.990 0.385 1.150 ;
  END
END BUFFD0

#--------EOF---------

MACRO BUFFD1
  CLASS CORE ;
  FOREIGN BUFFD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 2.045 1.410 2.305 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.780 0.800 4.600 ;
        RECT 0.585 2.480 0.885 2.780 ;
        RECT 0.670 1.280 0.800 2.480 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.710 0.815 3.190 ;
        RECT 0.605 2.550 0.865 2.710 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 1.065 2.085 1.760 2.215 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 2.230 0.335 4.970 ;
        RECT 0.175 2.070 1.345 2.230 ;
        RECT 0.175 1.150 0.335 2.070 ;
        RECT 0.125 0.990 0.385 1.150 ;
  END
END BUFFD1

#--------EOF---------

MACRO BUFFD2
  CLASS CORE ;
  FOREIGN BUFFD2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 0.670 2.085 1.845 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 1.615 1.570 1.775 2.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.615 1.410 3.265 1.570 ;
  END
END BUFFD2

#--------EOF---------

MACRO BUFFD4
  CLASS CORE ;
  FOREIGN BUFFD4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 3.005 1.410 5.185 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 0.585 2.085 1.760 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 2.025 2.085 5.600 2.215 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 2.230 1.295 4.070 ;
        RECT 1.135 2.070 2.305 2.230 ;
        RECT 1.135 1.570 1.295 2.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
  END
END BUFFD4

#--------EOF---------

MACRO BUFFD6
  CLASS CORE ;
  FOREIGN BUFFD6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 0.585 2.085 1.760 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.780800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 3.005 1.410 7.105 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 2.505 2.085 7.520 2.215 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 2.230 1.295 4.070 ;
        RECT 1.135 2.070 2.785 2.230 ;
        RECT 1.135 1.570 1.295 2.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
  END
END BUFFD6

#--------EOF---------

MACRO BUFFD8
  CLASS CORE ;
  FOREIGN BUFFD8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.220 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666900 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.395 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 0.585 2.085 2.720 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.405 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.374400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 7.805 4.070 8.065 4.230 ;
        RECT 9.725 4.070 9.985 4.230 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 7.855 1.570 8.015 4.070 ;
        RECT 9.775 1.570 9.935 4.070 ;
        RECT 3.965 1.410 9.985 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 11.220 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 11.220 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 3.465 2.085 10.400 2.215 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 2.230 2.255 4.070 ;
        RECT 2.095 2.070 3.745 2.230 ;
        RECT 2.095 1.570 2.255 2.070 ;
        RECT 0.125 1.410 2.305 1.570 ;
  END
END BUFFD8

#--------EOF---------

MACRO BUFFD12
  CLASS CORE ;
  FOREIGN BUFFD12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.000 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747500 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 0.670 4.215 0.800 4.480 ;
        RECT 1.630 4.215 1.760 4.480 ;
        RECT 2.590 4.215 2.720 4.480 ;
        RECT 3.550 4.215 3.680 4.480 ;
        RECT 4.510 4.215 4.640 4.480 ;
        RECT 0.670 4.085 4.640 4.215 ;
        RECT 0.670 2.300 0.800 4.085 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.555 0.800 2.000 ;
        RECT 0.670 1.425 4.640 1.555 ;
        RECT 0.670 1.350 0.800 1.425 ;
        RECT 1.630 1.350 1.760 1.425 ;
        RECT 2.590 1.350 2.720 1.425 ;
        RECT 3.550 1.350 3.680 1.425 ;
        RECT 4.510 1.350 4.640 1.425 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.561600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 7.805 4.070 8.065 4.230 ;
        RECT 9.725 4.070 9.985 4.230 ;
        RECT 11.645 4.070 11.905 4.230 ;
        RECT 13.565 4.070 13.825 4.230 ;
        RECT 15.485 4.070 15.745 4.230 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 7.855 1.570 8.015 4.070 ;
        RECT 9.775 1.570 9.935 4.070 ;
        RECT 11.695 1.570 11.855 4.070 ;
        RECT 13.615 1.570 13.775 4.070 ;
        RECT 15.535 1.570 15.695 4.070 ;
        RECT 5.885 1.410 15.745 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 16.445 0.990 16.705 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 12.655 0.150 12.815 0.990 ;
        RECT 14.575 0.150 14.735 0.990 ;
        RECT 16.495 0.150 16.655 0.990 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 17.000 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 12.655 5.130 12.815 5.970 ;
        RECT 14.575 5.130 14.735 5.970 ;
        RECT 16.495 5.130 16.655 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 14.525 4.970 14.785 5.130 ;
        RECT 16.445 4.970 16.705 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 16.030 5.200 16.160 5.380 ;
        RECT 5.470 2.300 5.600 4.000 ;
        RECT 5.385 2.215 5.685 2.300 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 14.110 2.215 14.240 4.000 ;
        RECT 15.070 2.215 15.200 4.000 ;
        RECT 16.030 2.215 16.160 4.000 ;
        RECT 5.385 2.085 16.160 2.215 ;
        RECT 5.385 2.000 5.685 2.085 ;
        RECT 5.470 1.640 5.600 2.000 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 14.110 1.640 14.240 2.085 ;
        RECT 15.070 1.640 15.200 2.085 ;
        RECT 16.030 1.640 16.160 2.085 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
        RECT 16.030 0.740 16.160 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 2.305 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 4.015 2.230 4.175 4.630 ;
        RECT 4.015 2.070 5.665 2.230 ;
        RECT 4.015 1.570 4.175 2.070 ;
        RECT 0.655 1.410 4.175 1.570 ;
        RECT 0.655 1.150 0.815 1.410 ;
        RECT 2.095 1.150 2.255 1.410 ;
        RECT 4.015 1.150 4.175 1.410 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
  END
END BUFFD12

#--------EOF---------

MACRO BUFFD16
  CLASS CORE ;
  FOREIGN BUFFD16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.331850 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 2.215 0.800 4.805 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 0.670 2.085 5.600 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 0.585 1.340 0.885 1.640 ;
        RECT 0.670 1.170 0.800 1.340 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 1.570 0.815 2.230 ;
        RECT 0.605 1.410 0.865 1.570 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.748799 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 10.685 4.070 10.945 4.230 ;
        RECT 12.605 4.070 12.865 4.230 ;
        RECT 14.525 4.070 14.785 4.230 ;
        RECT 16.445 4.070 16.705 4.230 ;
        RECT 18.365 4.070 18.625 4.230 ;
        RECT 20.285 4.070 20.545 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 8.815 1.570 8.975 4.070 ;
        RECT 10.735 1.570 10.895 4.070 ;
        RECT 12.655 1.570 12.815 4.070 ;
        RECT 14.575 1.570 14.735 4.070 ;
        RECT 16.495 1.570 16.655 4.070 ;
        RECT 18.415 1.570 18.575 4.070 ;
        RECT 20.335 1.570 20.495 4.070 ;
        RECT 6.845 1.410 20.545 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 15.485 0.990 15.745 1.150 ;
        RECT 17.405 0.990 17.665 1.150 ;
        RECT 19.325 0.990 19.585 1.150 ;
        RECT 21.245 0.990 21.505 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 15.535 0.150 15.695 0.990 ;
        RECT 17.455 0.150 17.615 0.990 ;
        RECT 19.375 0.150 19.535 0.990 ;
        RECT 21.295 0.150 21.455 0.990 ;
        RECT 0.000 -0.150 21.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 21.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 11.695 5.130 11.855 5.970 ;
        RECT 13.615 5.130 13.775 5.970 ;
        RECT 15.535 5.130 15.695 5.970 ;
        RECT 17.455 5.130 17.615 5.970 ;
        RECT 19.375 5.130 19.535 5.970 ;
        RECT 21.295 5.130 21.455 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
        RECT 13.565 4.970 13.825 5.130 ;
        RECT 15.485 4.970 15.745 5.130 ;
        RECT 17.405 4.970 17.665 5.130 ;
        RECT 19.325 4.970 19.585 5.130 ;
        RECT 21.245 4.970 21.505 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 16.030 5.200 16.160 5.380 ;
        RECT 16.990 5.200 17.120 5.380 ;
        RECT 17.950 5.200 18.080 5.380 ;
        RECT 18.910 5.200 19.040 5.380 ;
        RECT 19.870 5.200 20.000 5.380 ;
        RECT 20.830 5.200 20.960 5.380 ;
        RECT 6.430 2.300 6.560 4.000 ;
        RECT 6.345 2.215 6.645 2.300 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 14.110 2.215 14.240 4.000 ;
        RECT 15.070 2.215 15.200 4.000 ;
        RECT 16.030 2.215 16.160 4.000 ;
        RECT 16.990 2.215 17.120 4.000 ;
        RECT 17.950 2.215 18.080 4.000 ;
        RECT 18.910 2.215 19.040 4.000 ;
        RECT 19.870 2.215 20.000 4.000 ;
        RECT 20.830 2.215 20.960 4.000 ;
        RECT 6.345 2.085 20.960 2.215 ;
        RECT 6.345 2.000 6.645 2.085 ;
        RECT 6.430 1.640 6.560 2.000 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 14.110 1.640 14.240 2.085 ;
        RECT 15.070 1.640 15.200 2.085 ;
        RECT 16.030 1.640 16.160 2.085 ;
        RECT 16.990 1.640 17.120 2.085 ;
        RECT 17.950 1.640 18.080 2.085 ;
        RECT 18.910 1.640 19.040 2.085 ;
        RECT 19.870 1.640 20.000 2.085 ;
        RECT 20.830 1.640 20.960 2.085 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
        RECT 16.030 0.740 16.160 0.920 ;
        RECT 16.990 0.740 17.120 0.920 ;
        RECT 17.950 0.740 18.080 0.920 ;
        RECT 18.910 0.740 19.040 0.920 ;
        RECT 19.870 0.740 20.000 0.920 ;
        RECT 20.830 0.740 20.960 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 4.975 2.230 5.135 4.070 ;
        RECT 4.975 2.070 6.625 2.230 ;
        RECT 4.975 1.570 5.135 2.070 ;
        RECT 1.085 1.410 5.185 1.570 ;
  END
END BUFFD16

#--------EOF---------

MACRO DEL0
  CLASS CORE ;
  FOREIGN DEL0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 4.925 1.410 5.185 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 3.260 1.760 4.160 ;
        RECT 1.545 2.960 1.845 3.260 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 0.105 2.085 3.680 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 3.550 1.400 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.960 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 1.545 0.475 1.845 0.560 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 1.545 0.345 3.285 0.475 ;
        RECT 1.545 0.260 1.845 0.345 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 4.655 4.790 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 2.230 0.335 4.070 ;
        RECT 1.565 3.030 1.825 3.190 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 1.615 0.490 1.775 3.030 ;
        RECT 2.095 1.570 2.255 4.630 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 4.495 3.190 4.655 4.630 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END DEL0

#--------EOF---------

MACRO DEL01
  CLASS CORE ;
  FOREIGN DEL01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 4.925 1.410 5.185 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 3.260 1.760 4.000 ;
        RECT 1.545 3.175 1.845 3.260 ;
        RECT 2.985 3.175 3.285 3.260 ;
        RECT 1.545 3.045 3.285 3.175 ;
        RECT 1.545 2.960 1.845 3.045 ;
        RECT 2.985 2.960 3.285 3.045 ;
        RECT 0.105 2.695 0.405 2.780 ;
        RECT 3.550 2.695 3.680 4.000 ;
        RECT 0.105 2.565 3.680 2.695 ;
        RECT 0.105 2.480 0.405 2.565 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 0.105 2.085 3.680 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 4.000 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 1.545 0.260 1.845 0.560 ;
        RECT 2.025 0.475 2.325 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 2.025 0.345 4.640 0.475 ;
        RECT 2.025 0.260 2.325 0.345 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 0.175 2.710 0.335 4.070 ;
        RECT 1.565 3.030 1.825 3.190 ;
        RECT 0.125 2.550 0.385 2.710 ;
        RECT 0.175 2.230 0.335 2.550 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 1.615 1.150 1.775 3.030 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 3.055 3.190 3.215 4.070 ;
        RECT 3.005 3.030 3.265 3.190 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 1.615 0.990 3.265 1.150 ;
        RECT 1.615 0.490 1.775 0.990 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 2.045 0.330 2.305 0.490 ;
  END
END DEL01

#--------EOF---------

MACRO DEL02
  CLASS CORE ;
  FOREIGN DEL02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 6.845 1.410 7.105 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 1.630 2.215 1.760 4.635 ;
        RECT 0.105 2.085 1.760 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.255 1.760 2.085 ;
        RECT 2.590 1.255 2.720 4.635 ;
        RECT 4.510 4.215 4.640 4.635 ;
        RECT 5.470 4.215 5.600 4.635 ;
        RECT 4.510 4.085 5.600 4.215 ;
        RECT 4.510 1.255 4.640 1.435 ;
        RECT 5.470 1.255 5.600 4.085 ;
        RECT 5.865 3.175 6.165 3.260 ;
        RECT 7.390 3.175 7.520 4.000 ;
        RECT 5.865 3.045 7.520 3.175 ;
        RECT 5.865 2.960 6.165 3.045 ;
        RECT 5.865 2.215 6.165 2.300 ;
        RECT 5.865 2.085 7.520 2.215 ;
        RECT 5.865 2.000 6.165 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 1.630 0.345 2.720 0.475 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 2.985 0.345 5.600 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 2.230 0.335 4.070 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 2.095 1.150 2.255 4.970 ;
        RECT 3.055 1.150 3.215 4.970 ;
        RECT 4.975 1.150 5.135 4.970 ;
        RECT 5.935 3.190 6.095 4.970 ;
        RECT 5.885 3.030 6.145 3.190 ;
        RECT 5.935 2.230 6.095 3.030 ;
        RECT 5.885 2.070 6.145 2.230 ;
        RECT 5.935 1.150 6.095 2.070 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END DEL02

#--------EOF---------

MACRO DEL2
  CLASS CORE ;
  FOREIGN DEL2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 4.925 1.410 5.185 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 4.215 1.760 4.300 ;
        RECT 2.505 4.215 2.805 4.300 ;
        RECT 1.630 4.085 2.805 4.215 ;
        RECT 2.505 4.000 2.805 4.085 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 0.105 2.085 3.680 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 3.550 1.400 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.960 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 1.630 0.345 3.285 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 4.655 4.790 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 2.230 0.335 4.070 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 2.095 1.570 2.255 4.630 ;
        RECT 2.525 4.070 3.265 4.230 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 4.495 3.190 4.655 4.630 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END DEL2

#--------EOF---------

MACRO DEL4
  CLASS CORE ;
  FOREIGN DEL4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 4.925 1.410 5.185 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 4.215 1.760 4.350 ;
        RECT 2.505 4.215 2.805 4.300 ;
        RECT 1.630 4.085 2.805 4.215 ;
        RECT 2.505 4.000 2.805 4.085 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 0.105 2.085 3.680 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 3.550 1.400 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.960 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 1.630 0.345 3.285 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 4.655 4.790 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 2.230 0.335 4.070 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 2.095 1.570 2.255 4.630 ;
        RECT 2.525 4.070 3.265 4.230 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 4.495 3.190 4.655 4.630 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END DEL4

#--------EOF---------

MACRO DEL005
  CLASS CORE ;
  FOREIGN DEL005 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.422500 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 0.670 3.045 1.760 3.175 ;
        RECT 0.670 1.345 0.800 3.045 ;
        RECT 1.630 1.345 1.760 1.525 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 0.585 0.345 1.760 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
      LAYER Metal1 ;
        RECT 0.655 0.490 0.815 1.150 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 3.005 1.410 3.265 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 3.260 2.720 4.000 ;
        RECT 2.505 2.960 2.805 3.260 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 1.065 2.085 2.720 2.215 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 3.190 0.335 4.070 ;
        RECT 0.175 3.030 2.785 3.190 ;
        RECT 0.175 2.230 0.335 3.030 ;
        RECT 0.175 2.070 1.345 2.230 ;
        RECT 0.175 1.150 0.335 2.070 ;
        RECT 0.125 0.990 0.385 1.150 ;
  END
END DEL005

#--------EOF---------

MACRO DEL015
  CLASS CORE ;
  FOREIGN DEL015 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 6.845 1.410 7.105 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.260 0.800 4.000 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.030 0.865 3.190 ;
        RECT 0.655 0.490 0.815 3.030 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 0.105 2.085 1.760 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 4.000 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 4.510 1.640 4.640 3.045 ;
        RECT 5.470 1.640 5.600 1.820 ;
        RECT 7.390 1.640 7.520 4.000 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 1.630 0.345 2.720 0.475 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 7.390 0.560 7.520 0.920 ;
        RECT 2.985 0.345 5.600 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
        RECT 7.305 0.260 7.605 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 0.175 2.230 0.335 4.070 ;
        RECT 0.125 2.070 0.385 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 4.925 1.410 5.185 1.570 ;
        RECT 5.885 1.410 6.145 1.570 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 5.935 0.490 6.095 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 5.935 0.330 7.585 0.490 ;
  END
END DEL015

#--------EOF---------

MACRO DFCNQD1
  CLASS BLOCK ;
  FOREIGN DFCNQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.000 BY 6.120 ;
  SYMMETRY X Y R90 ;
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.155 0.800 4.650 ;
        RECT 0.190 3.025 0.800 3.155 ;
        RECT 0.190 2.280 0.320 3.025 ;
        RECT 0.105 1.980 0.405 2.280 ;
        RECT 0.190 1.535 0.320 1.980 ;
        RECT 0.190 1.405 0.800 1.535 ;
        RECT 0.670 1.270 0.800 1.405 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 2.210 0.335 2.690 ;
        RECT 0.125 2.050 0.385 2.210 ;
    END
  END cp
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150800 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.390 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.270 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 1.390 4.655 2.050 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.287300 ;
    PORT
      LAYER GatPoly ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 8.350 4.775 8.480 4.925 ;
        RECT 7.390 4.645 8.480 4.775 ;
        RECT 7.390 1.940 7.520 4.645 ;
        RECT 13.150 3.720 13.280 4.210 ;
        RECT 13.065 3.420 13.365 3.720 ;
        RECT 13.065 1.980 13.365 2.280 ;
        RECT 7.305 1.640 7.605 1.940 ;
        RECT 7.390 1.165 7.520 1.640 ;
        RECT 13.150 1.620 13.280 1.980 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
      LAYER Metal1 ;
        RECT 13.085 3.490 13.345 3.650 ;
        RECT 13.135 2.210 13.295 3.490 ;
        RECT 11.215 2.050 13.345 2.210 ;
        RECT 11.215 1.870 11.375 2.050 ;
        RECT 7.325 1.710 11.375 1.870 ;
    END
  END cdn
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.485 4.630 16.655 4.790 ;
        RECT 16.495 1.150 16.655 4.630 ;
        RECT 16.445 0.990 16.705 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 12.605 0.990 15.745 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.005 0.650 3.265 0.810 ;
        RECT 3.055 0.150 3.215 0.650 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 15.535 0.150 15.695 0.990 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 17.000 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 6.895 5.470 7.055 5.970 ;
        RECT 8.815 5.470 8.975 5.970 ;
        RECT 12.655 5.470 12.815 5.970 ;
        RECT 6.845 5.310 7.105 5.470 ;
        RECT 8.765 5.310 9.025 5.470 ;
        RECT 12.605 5.310 12.865 5.470 ;
        RECT 14.575 5.130 14.735 5.970 ;
        RECT 1.085 4.970 3.265 5.130 ;
        RECT 14.525 4.970 14.785 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 5.385 5.560 5.685 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.560 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 5.470 4.690 5.600 4.870 ;
        RECT 1.630 2.760 1.760 4.650 ;
        RECT 3.550 3.720 3.680 4.390 ;
        RECT 6.430 3.720 6.560 4.895 ;
        RECT 3.465 3.420 3.765 3.720 ;
        RECT 6.345 3.420 6.645 3.720 ;
        RECT 0.585 2.675 0.885 2.760 ;
        RECT 1.545 2.675 1.845 2.760 ;
        RECT 0.585 2.545 1.845 2.675 ;
        RECT 0.585 2.460 0.885 2.545 ;
        RECT 1.545 2.460 1.845 2.545 ;
        RECT 1.630 1.270 1.760 2.460 ;
        RECT 3.550 2.280 3.680 3.420 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 6.430 1.940 6.560 3.420 ;
        RECT 8.265 2.940 8.565 3.240 ;
        RECT 8.350 2.280 8.480 2.940 ;
        RECT 9.310 2.280 9.440 4.485 ;
        RECT 10.270 2.760 10.400 4.170 ;
        RECT 10.185 2.460 10.485 2.760 ;
        RECT 8.265 1.980 8.565 2.280 ;
        RECT 9.225 1.980 9.525 2.280 ;
        RECT 6.345 1.640 6.645 1.940 ;
        RECT 2.505 1.535 2.805 1.620 ;
        RECT 2.505 1.405 3.680 1.535 ;
        RECT 2.505 1.320 2.805 1.405 ;
        RECT 3.550 1.270 3.680 1.405 ;
        RECT 5.470 1.165 5.600 1.345 ;
        RECT 6.430 1.165 6.560 1.640 ;
        RECT 8.350 1.350 8.480 1.980 ;
        RECT 9.310 1.410 9.440 1.590 ;
        RECT 10.270 1.165 10.400 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 5.470 0.560 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 5.385 0.475 5.685 0.560 ;
        RECT 9.310 0.475 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.475 11.360 4.925 ;
        RECT 12.190 3.155 12.320 4.925 ;
        RECT 14.110 3.720 14.240 4.210 ;
        RECT 14.025 3.420 14.325 3.720 ;
        RECT 13.545 3.155 13.845 3.240 ;
        RECT 15.070 3.155 15.200 4.100 ;
        RECT 12.190 3.025 16.160 3.155 ;
        RECT 12.190 1.620 12.320 3.025 ;
        RECT 13.545 2.940 13.845 3.025 ;
        RECT 14.025 2.460 14.325 2.760 ;
        RECT 14.110 1.620 14.240 2.460 ;
        RECT 16.030 1.620 16.160 3.025 ;
        RECT 12.105 1.320 12.405 1.620 ;
        RECT 12.190 1.165 12.320 1.320 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 14.110 0.560 14.240 0.920 ;
        RECT 16.030 0.740 16.160 0.920 ;
        RECT 5.385 0.345 11.360 0.475 ;
        RECT 5.385 0.260 5.685 0.345 ;
        RECT 14.025 0.260 14.325 0.560 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 5.665 5.790 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 5.885 4.970 8.065 5.130 ;
        RECT 10.685 4.970 14.255 5.130 ;
        RECT 0.655 2.690 0.815 4.970 ;
        RECT 2.045 4.610 3.695 4.770 ;
        RECT 4.925 4.630 5.615 4.790 ;
        RECT 3.535 3.650 3.695 4.610 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 5.455 3.170 5.615 4.630 ;
        RECT 9.295 4.630 9.985 4.790 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 9.295 3.650 9.455 4.630 ;
        RECT 6.365 3.490 9.455 3.650 ;
        RECT 13.615 3.170 13.775 4.630 ;
        RECT 14.095 3.650 14.255 4.970 ;
        RECT 14.045 3.490 14.305 3.650 ;
        RECT 5.455 3.010 8.545 3.170 ;
        RECT 13.565 3.010 13.825 3.170 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 2.575 2.530 10.465 2.690 ;
        RECT 1.615 1.550 1.775 2.530 ;
        RECT 2.575 1.550 2.735 2.530 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 4.975 2.050 9.505 2.210 ;
        RECT 0.175 1.390 2.785 1.550 ;
        RECT 0.175 1.150 0.335 1.390 ;
        RECT 3.535 1.150 3.695 2.050 ;
        RECT 4.975 1.150 5.135 2.050 ;
        RECT 6.365 1.710 6.625 1.870 ;
        RECT 6.415 1.530 6.575 1.710 ;
        RECT 13.615 1.550 13.775 3.010 ;
        RECT 14.095 2.690 14.255 3.490 ;
        RECT 14.045 2.530 14.305 2.690 ;
        RECT 6.415 1.370 8.975 1.530 ;
        RECT 12.125 1.390 14.785 1.550 ;
        RECT 8.815 1.150 8.975 1.370 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 3.695 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 10.685 0.990 11.905 1.150 ;
        RECT 3.535 0.490 3.695 0.990 ;
        RECT 9.775 0.490 9.935 0.990 ;
        RECT 3.535 0.330 5.665 0.490 ;
        RECT 9.775 0.330 14.305 0.490 ;
  END
END DFCNQD1

#--------EOF---------

MACRO DFQD1
  CLASS CORE ;
  FOREIGN DFQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.152100 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 4.215 4.640 4.450 ;
        RECT 4.905 4.215 5.205 4.300 ;
        RECT 4.510 4.085 5.205 4.215 ;
        RECT 4.905 4.000 5.205 4.085 ;
        RECT 4.990 2.695 5.120 4.000 ;
        RECT 4.510 2.565 5.120 2.695 ;
        RECT 4.510 1.340 4.640 2.565 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.975 4.230 5.135 4.790 ;
        RECT 4.925 4.070 5.185 4.230 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.780 1.760 4.000 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 1.640 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.550 2.255 2.710 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 12.605 4.070 12.865 4.230 ;
        RECT 12.655 1.570 12.815 4.070 ;
        RECT 12.605 1.410 12.865 1.570 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 13.615 5.130 13.775 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 13.565 4.970 13.825 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.025 5.775 2.325 5.860 ;
        RECT 5.865 5.775 6.165 5.860 ;
        RECT 0.670 5.645 5.600 5.775 ;
        RECT 0.670 5.200 0.800 5.645 ;
        RECT 2.025 5.560 2.325 5.645 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 5.865 5.645 7.520 5.775 ;
        RECT 5.865 5.560 6.165 5.645 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.645 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 5.470 4.720 5.600 4.900 ;
        RECT 2.505 4.000 2.805 4.300 ;
        RECT 0.670 1.640 0.800 4.000 ;
        RECT 2.590 1.220 2.720 4.000 ;
        RECT 3.550 3.260 3.680 4.315 ;
        RECT 6.430 4.300 6.560 4.900 ;
        RECT 6.345 4.000 6.645 4.300 ;
        RECT 3.465 2.960 3.765 3.260 ;
        RECT 5.385 2.960 5.685 3.260 ;
        RECT 3.465 2.480 3.765 2.780 ;
        RECT 3.550 1.340 3.680 2.480 ;
        RECT 2.505 0.920 2.805 1.220 ;
        RECT 5.470 1.170 5.600 2.960 ;
        RECT 6.430 1.640 6.560 4.000 ;
        RECT 6.345 1.340 6.645 1.640 ;
        RECT 7.390 1.390 7.520 4.450 ;
        RECT 8.350 2.780 8.480 4.135 ;
        RECT 9.310 3.260 9.440 4.900 ;
        RECT 9.225 2.960 9.525 3.260 ;
        RECT 8.265 2.695 8.565 2.780 ;
        RECT 8.265 2.565 8.960 2.695 ;
        RECT 8.265 2.480 8.565 2.565 ;
        RECT 8.265 2.000 8.565 2.300 ;
        RECT 6.430 1.170 6.560 1.340 ;
        RECT 8.350 1.305 8.480 2.000 ;
        RECT 8.830 1.555 8.960 2.565 ;
        RECT 10.270 2.300 10.400 4.900 ;
        RECT 10.185 2.000 10.485 2.300 ;
        RECT 8.830 1.425 9.440 1.555 ;
        RECT 9.310 1.170 9.440 1.425 ;
        RECT 10.270 1.170 10.400 2.000 ;
        RECT 11.230 1.640 11.360 4.000 ;
        RECT 11.625 2.215 11.925 2.300 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 11.625 2.085 13.280 2.215 ;
        RECT 11.625 2.000 11.925 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 0.670 0.345 3.680 0.475 ;
        RECT 4.905 0.475 5.205 0.560 ;
        RECT 7.390 0.475 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 4.905 0.345 7.520 0.475 ;
        RECT 8.745 0.475 9.045 0.560 ;
        RECT 9.705 0.475 10.005 0.560 ;
        RECT 11.230 0.475 11.360 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 8.745 0.345 11.360 0.475 ;
        RECT 4.905 0.260 5.205 0.345 ;
        RECT 8.745 0.260 9.045 0.345 ;
        RECT 9.705 0.260 10.005 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 5.630 2.305 5.790 ;
        RECT 4.975 5.630 6.145 5.790 ;
        RECT 2.095 5.130 2.255 5.630 ;
        RECT 4.975 5.130 5.135 5.630 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 7.855 4.230 8.015 4.630 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.785 4.230 ;
        RECT 6.365 4.070 8.015 4.230 ;
        RECT 8.815 4.230 8.975 4.630 ;
        RECT 8.815 4.070 9.935 4.230 ;
        RECT 11.645 4.070 11.905 4.230 ;
        RECT 0.175 3.190 0.335 4.070 ;
        RECT 0.175 3.030 9.505 3.190 ;
        RECT 3.485 2.550 8.545 2.710 ;
        RECT 8.815 2.230 8.975 3.030 ;
        RECT 0.175 2.070 8.975 2.230 ;
        RECT 0.175 1.570 0.335 2.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
        RECT 6.365 1.410 8.015 1.570 ;
        RECT 7.855 1.150 8.015 1.410 ;
        RECT 2.045 0.990 2.785 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 8.815 0.490 8.975 0.990 ;
        RECT 9.775 0.490 9.935 4.070 ;
        RECT 11.695 2.230 11.855 4.070 ;
        RECT 10.205 2.070 11.905 2.230 ;
        RECT 11.695 1.570 11.855 2.070 ;
        RECT 11.645 1.410 11.905 1.570 ;
        RECT 4.925 0.330 5.185 0.490 ;
        RECT 8.765 0.330 9.025 0.490 ;
        RECT 9.725 0.330 9.985 0.490 ;
  END
END DFQD1

#--------EOF---------

MACRO FILL1
  CLASS CORE ;
  FOREIGN FILL1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.340 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.340 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 0.340 6.270 ;
    END
  END vdd
END FILL1

#--------EOF---------

MACRO FILL2
  CLASS CORE ;
  FOREIGN FILL2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.680 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.680 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 0.680 6.270 ;
    END
  END vdd
END FILL2

#--------EOF---------

MACRO FILL4
  CLASS CORE ;
  FOREIGN FILL4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.360 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 1.360 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.360 6.270 ;
    END
  END vdd
END FILL4

#--------EOF---------

MACRO FILL8
  CLASS CORE ;
  FOREIGN FILL8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END FILL8

#--------EOF---------

MACRO INVD0
  CLASS CORE ;
  FOREIGN INVD0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
    END
  END vdd
END INVD0

#--------EOF---------

MACRO INVD1
  CLASS CORE ;
  FOREIGN INVD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
END INVD1

#--------EOF---------

MACRO INVD2
  CLASS CORE ;
  FOREIGN INVD2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 0.670 2.085 1.845 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
END INVD2

#--------EOF---------

MACRO INVD4
  CLASS CORE ;
  FOREIGN INVD4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.085 1.410 3.265 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 0.670 2.085 3.765 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
END INVD4

#--------EOF---------

MACRO INVD6
  CLASS CORE ;
  FOREIGN INVD6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.356800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 0.125 1.410 6.145 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.497600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 0.585 2.085 5.600 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
END INVD6

#--------EOF---------

MACRO INVD8
  CLASS CORE ;
  FOREIGN INVD8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.950400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 7.805 4.070 8.065 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 7.855 1.570 8.015 4.070 ;
        RECT 0.125 1.410 8.065 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.996800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 0.585 2.085 7.520 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
END INVD8

#--------EOF---------

MACRO INVD12
  CLASS CORE ;
  FOREIGN INVD12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.137600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 7.805 4.070 8.065 4.230 ;
        RECT 9.725 4.070 9.985 4.230 ;
        RECT 11.645 4.070 11.905 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 7.855 1.570 8.015 4.070 ;
        RECT 9.775 1.570 9.935 4.070 ;
        RECT 11.695 1.570 11.855 4.070 ;
        RECT 0.125 1.410 11.905 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.995200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 0.585 2.085 11.360 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
    END
  END vdd
END INVD12

#--------EOF---------

MACRO INVD16
  CLASS CORE ;
  FOREIGN INVD16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.980 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.324800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 7.805 4.070 8.065 4.230 ;
        RECT 9.725 4.070 9.985 4.230 ;
        RECT 11.645 4.070 11.905 4.230 ;
        RECT 13.565 4.070 13.825 4.230 ;
        RECT 15.485 4.070 15.745 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 7.855 1.570 8.015 4.070 ;
        RECT 9.775 1.570 9.935 4.070 ;
        RECT 11.695 1.570 11.855 4.070 ;
        RECT 13.615 1.570 13.775 4.070 ;
        RECT 15.535 1.570 15.695 4.070 ;
        RECT 0.125 1.410 15.745 1.570 ;
    END
  END zn
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.993600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 8.350 2.215 8.480 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 14.110 2.215 14.240 4.000 ;
        RECT 15.070 2.215 15.200 4.000 ;
        RECT 0.585 2.085 15.200 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 8.350 1.640 8.480 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 14.110 1.640 14.240 2.085 ;
        RECT 15.070 1.640 15.200 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 12.655 0.150 12.815 0.990 ;
        RECT 14.575 0.150 14.735 0.990 ;
        RECT 0.000 -0.150 15.980 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 15.980 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 12.655 5.130 12.815 5.970 ;
        RECT 14.575 5.130 14.735 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 14.525 4.970 14.785 5.130 ;
    END
  END vdd
END INVD16

#--------EOF---------

MACRO MUX2D0
  CLASS CORE ;
  FOREIGN MUX2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 4.215 2.720 4.600 ;
        RECT 4.510 4.215 4.640 4.600 ;
        RECT 1.150 4.085 4.640 4.215 ;
        RECT 1.150 2.215 1.280 4.085 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 1.150 2.085 1.845 2.215 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 4.510 1.280 4.640 4.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 1.615 1.410 1.775 2.070 ;
    END
  END s
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 3.465 5.560 3.765 5.860 ;
        RECT 3.550 5.200 3.680 5.560 ;
        RECT 3.550 4.420 3.680 4.600 ;
        RECT 3.465 2.960 3.765 3.260 ;
        RECT 3.550 1.280 3.680 2.960 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 3.535 3.190 3.695 5.630 ;
        RECT 3.485 3.030 3.745 3.190 ;
    END
  END i0
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 1.150 6.095 4.970 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 4.420 1.760 4.600 ;
        RECT 1.545 2.695 1.845 2.780 ;
        RECT 2.985 2.695 3.285 2.780 ;
        RECT 1.545 2.565 3.285 2.695 ;
        RECT 1.545 2.480 1.845 2.565 ;
        RECT 2.590 1.280 2.720 2.565 ;
        RECT 2.985 2.480 3.285 2.565 ;
        RECT 6.430 1.280 6.560 4.600 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 2.025 0.475 2.325 0.560 ;
        RECT 6.430 0.475 6.560 0.920 ;
        RECT 2.025 0.345 6.560 0.475 ;
        RECT 2.025 0.260 2.325 0.345 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 1.615 2.710 1.775 5.630 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.575 4.970 3.265 5.130 ;
        RECT 4.495 4.970 5.185 5.130 ;
        RECT 1.565 2.550 1.825 2.710 ;
        RECT 2.095 1.150 2.255 4.970 ;
        RECT 2.575 1.150 2.735 4.970 ;
        RECT 4.495 2.710 4.655 4.970 ;
        RECT 3.005 2.550 5.135 2.710 ;
        RECT 4.975 1.150 5.135 2.550 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.575 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 2.045 0.330 2.305 0.490 ;
  END
END MUX2D0

#--------EOF---------

MACRO MUX2D1
  CLASS CORE ;
  FOREIGN MUX2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.545 5.775 1.845 5.860 ;
        RECT 1.545 5.645 4.640 5.775 ;
        RECT 1.545 5.560 1.845 5.645 ;
        RECT 2.590 5.200 2.720 5.645 ;
        RECT 4.510 5.200 4.640 5.645 ;
        RECT 2.590 4.420 2.720 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 4.510 1.280 4.640 4.600 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 1.615 2.230 1.775 5.630 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196300 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.780 3.680 4.210 ;
        RECT 3.465 2.480 3.765 2.780 ;
        RECT 3.550 1.440 3.680 2.480 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.710 3.695 3.190 ;
        RECT 3.485 2.550 3.745 2.710 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.881400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.570 6.095 4.630 ;
        RECT 5.885 1.410 6.145 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 4.215 1.760 4.600 ;
        RECT 1.630 4.085 2.720 4.215 ;
        RECT 2.590 2.215 2.720 4.085 ;
        RECT 2.985 2.215 3.285 2.300 ;
        RECT 2.590 2.085 3.285 2.215 ;
        RECT 2.590 1.280 2.720 2.085 ;
        RECT 2.985 2.000 3.285 2.085 ;
        RECT 6.430 1.640 6.560 4.360 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 2.025 0.475 2.325 0.560 ;
        RECT 6.430 0.475 6.560 0.920 ;
        RECT 2.025 0.345 6.560 0.475 ;
        RECT 2.025 0.260 2.325 0.345 ;
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
        RECT 2.095 1.150 2.255 4.970 ;
        RECT 2.575 4.630 3.265 4.790 ;
        RECT 2.575 1.150 2.735 4.630 ;
        RECT 4.975 2.230 5.135 4.970 ;
        RECT 3.005 2.070 5.135 2.230 ;
        RECT 4.975 1.150 5.135 2.070 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.575 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 2.045 0.330 2.305 0.490 ;
  END
END MUX2D1

#--------EOF---------

MACRO MUX2D2
  CLASS CORE ;
  FOREIGN MUX2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.505 5.560 2.805 5.860 ;
        RECT 2.590 5.200 2.720 5.560 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 4.420 2.720 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 4.510 1.280 4.640 4.600 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 1.630 0.345 4.640 0.475 ;
      LAYER Metal1 ;
        RECT 1.615 5.630 2.785 5.790 ;
        RECT 1.615 2.230 1.775 5.630 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196300 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.210 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.440 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 6.845 1.410 7.105 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.985 5.775 3.285 5.860 ;
        RECT 2.985 5.645 6.560 5.775 ;
        RECT 2.985 5.560 3.285 5.645 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 6.430 5.200 6.560 5.645 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 1.630 4.215 1.760 4.600 ;
        RECT 1.630 4.085 2.720 4.215 ;
        RECT 2.590 3.175 2.720 4.085 ;
        RECT 2.985 3.175 3.285 3.260 ;
        RECT 2.590 3.045 3.285 3.175 ;
        RECT 2.590 1.280 2.720 3.045 ;
        RECT 2.985 2.960 3.285 3.045 ;
        RECT 6.430 3.175 6.560 4.000 ;
        RECT 7.390 3.175 7.520 4.000 ;
        RECT 6.430 3.045 7.520 3.175 ;
        RECT 6.430 1.640 6.560 3.045 ;
        RECT 7.390 1.640 7.520 1.820 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 6.430 0.475 6.560 0.920 ;
        RECT 7.390 0.475 7.520 0.920 ;
        RECT 6.430 0.345 7.520 0.475 ;
      LAYER Metal1 ;
        RECT 3.005 5.630 3.265 5.790 ;
        RECT 3.055 5.130 3.215 5.630 ;
        RECT 2.045 4.970 3.215 5.130 ;
        RECT 4.495 4.970 5.185 5.130 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
        RECT 2.095 1.150 2.255 4.970 ;
        RECT 2.575 4.630 3.265 4.790 ;
        RECT 2.575 1.150 2.735 4.630 ;
        RECT 4.495 3.190 4.655 4.970 ;
        RECT 3.005 3.030 5.135 3.190 ;
        RECT 4.975 1.150 5.135 3.030 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.575 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
  END
END MUX2D2

#--------EOF---------

MACRO MUX2D4
  CLASS CORE ;
  FOREIGN MUX2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.347750 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 7.520 5.775 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 7.390 5.200 7.520 5.645 ;
        RECT 7.390 4.300 7.520 4.600 ;
        RECT 3.550 3.260 3.680 4.105 ;
        RECT 7.305 4.000 7.605 4.300 ;
        RECT 3.465 2.960 3.765 3.260 ;
        RECT 7.305 2.000 7.605 2.300 ;
        RECT 2.590 1.540 2.720 1.720 ;
        RECT 7.390 1.280 7.520 2.000 ;
        RECT 2.590 0.560 2.720 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 2.505 0.260 2.805 0.560 ;
      LAYER Metal1 ;
        RECT 7.325 4.070 7.585 4.230 ;
        RECT 3.485 3.030 3.745 3.190 ;
        RECT 3.535 0.490 3.695 3.030 ;
        RECT 7.375 2.230 7.535 4.070 ;
        RECT 7.325 2.070 7.585 2.230 ;
        RECT 2.525 0.330 3.695 0.490 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 0.670 3.045 1.760 3.175 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 1.630 1.640 1.760 3.045 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 0.585 0.345 1.760 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
      LAYER Metal1 ;
        RECT 0.655 0.490 0.815 1.150 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388700 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 4.510 3.175 4.640 4.225 ;
        RECT 5.470 3.260 5.600 4.225 ;
        RECT 5.385 3.175 5.685 3.260 ;
        RECT 4.510 3.045 5.685 3.175 ;
        RECT 5.385 2.960 5.685 3.045 ;
        RECT 5.385 2.215 5.685 2.300 ;
        RECT 4.510 2.085 5.685 2.215 ;
        RECT 4.510 1.440 4.640 2.085 ;
        RECT 5.385 2.000 5.685 2.085 ;
        RECT 5.470 1.440 5.600 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 5.405 3.030 5.665 3.190 ;
        RECT 5.455 2.230 5.615 3.030 ;
        RECT 5.405 2.070 5.665 2.230 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 10.685 4.070 10.945 4.230 ;
        RECT 8.815 1.570 8.975 4.070 ;
        RECT 10.735 1.570 10.895 4.070 ;
        RECT 8.765 1.410 10.945 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 11.695 5.130 11.855 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 8.350 3.175 8.480 4.000 ;
        RECT 9.310 3.175 9.440 4.000 ;
        RECT 10.270 3.175 10.400 4.000 ;
        RECT 11.230 3.175 11.360 4.000 ;
        RECT 8.350 3.045 11.360 3.175 ;
        RECT 2.985 2.695 3.285 2.780 ;
        RECT 9.310 2.695 9.440 3.045 ;
        RECT 2.985 2.565 9.440 2.695 ;
        RECT 2.985 2.480 3.285 2.565 ;
        RECT 2.590 2.085 3.680 2.215 ;
        RECT 3.550 1.455 3.680 2.085 ;
        RECT 8.350 1.640 8.480 1.820 ;
        RECT 9.310 1.640 9.440 2.565 ;
        RECT 10.270 1.640 10.400 3.045 ;
        RECT 11.230 1.640 11.360 1.820 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 6.825 0.475 7.125 0.560 ;
        RECT 3.550 0.345 7.125 0.475 ;
        RECT 8.350 0.475 8.480 0.920 ;
        RECT 9.310 0.475 9.440 0.920 ;
        RECT 10.270 0.475 10.400 0.920 ;
        RECT 11.230 0.475 11.360 0.920 ;
        RECT 8.350 0.345 11.360 0.475 ;
        RECT 6.825 0.260 7.125 0.345 ;
      LAYER Metal1 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 3.965 4.630 6.145 4.790 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 1.615 4.070 2.305 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 1.615 1.570 1.775 4.070 ;
        RECT 3.055 2.710 3.215 4.070 ;
        RECT 3.005 2.550 3.265 2.710 ;
        RECT 0.125 1.410 2.305 1.570 ;
        RECT 0.175 1.150 0.335 1.410 ;
        RECT 3.055 1.150 3.215 2.550 ;
        RECT 4.015 1.570 4.175 4.630 ;
        RECT 4.015 1.410 6.095 1.570 ;
        RECT 4.015 1.150 4.175 1.410 ;
        RECT 5.935 1.150 6.095 1.410 ;
        RECT 6.895 1.150 7.055 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.895 0.490 7.055 0.990 ;
        RECT 6.845 0.330 7.105 0.490 ;
  END
END MUX2D4

#--------EOF---------

MACRO ND2D0
  CLASS CORE ;
  FOREIGN ND2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.701400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 1.135 4.630 2.255 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
END ND2D0

#--------EOF---------

MACRO ND2D1
  CLASS CORE ;
  FOREIGN ND2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.402800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 3.190 1.295 4.070 ;
        RECT 1.135 3.030 2.255 3.190 ;
        RECT 2.095 1.570 2.255 3.030 ;
        RECT 2.045 1.410 2.305 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
END ND2D1

#--------EOF---------

MACRO ND2D2
  CLASS CORE ;
  FOREIGN ND2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.589600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.135 3.190 1.295 4.070 ;
        RECT 3.055 3.190 3.215 4.070 ;
        RECT 1.135 3.030 3.215 3.190 ;
        RECT 2.095 1.570 2.255 3.030 ;
        RECT 2.045 1.410 2.305 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 1.630 2.085 2.805 2.215 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 0.670 2.085 1.365 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 2.070 1.775 2.230 ;
        RECT 3.485 2.070 3.745 2.230 ;
        RECT 1.615 1.150 1.775 2.070 ;
        RECT 3.535 1.150 3.695 2.070 ;
        RECT 1.615 0.990 3.695 1.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
END ND2D2

#--------EOF---------

MACRO ND2D4
  CLASS CORE ;
  FOREIGN ND2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.179200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 3.265 4.230 ;
        RECT 4.925 4.070 7.105 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 4.975 1.570 5.135 4.070 ;
        RECT 2.045 1.410 6.145 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 1.630 2.085 6.560 2.215 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.670 1.640 0.800 4.000 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 5.470 3.260 5.600 4.000 ;
        RECT 5.385 3.175 5.685 3.260 ;
        RECT 4.510 3.045 5.685 3.175 ;
        RECT 5.385 2.960 5.685 3.045 ;
        RECT 6.825 3.175 7.125 3.260 ;
        RECT 7.390 3.175 7.520 4.000 ;
        RECT 6.825 3.045 7.520 3.175 ;
        RECT 6.825 2.960 7.125 3.045 ;
        RECT 6.910 2.215 7.040 2.960 ;
        RECT 6.910 2.085 7.520 2.215 ;
        RECT 3.550 1.640 3.680 1.820 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 7.390 0.475 7.520 0.920 ;
        RECT 0.670 0.345 7.520 0.475 ;
      LAYER Metal1 ;
        RECT 5.405 3.030 7.105 3.190 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
END ND2D4

#--------EOF---------

MACRO ND3D0
  CLASS CORE ;
  FOREIGN ND3D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.040400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 0.175 3.190 0.335 4.970 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 1.135 4.630 2.255 4.790 ;
        RECT 1.135 3.190 1.295 4.630 ;
        RECT 0.175 3.030 1.295 3.190 ;
        RECT 0.175 1.150 0.335 3.030 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
END ND3D0

#--------EOF---------

MACRO ND3D1
  CLASS CORE ;
  FOREIGN ND3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.815 4.230 ;
        RECT 0.655 2.710 0.815 4.070 ;
        RECT 1.615 4.070 2.305 4.230 ;
        RECT 1.615 2.710 1.775 4.070 ;
        RECT 0.655 2.550 1.775 2.710 ;
        RECT 0.655 1.570 0.815 2.550 ;
        RECT 0.125 1.410 0.815 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.105 2.215 0.405 2.300 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 0.105 2.085 0.800 2.215 ;
        RECT 0.105 2.000 0.405 2.085 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 2.230 0.335 2.710 ;
        RECT 0.125 2.070 0.385 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 1.615 1.410 1.775 2.070 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
END ND3D1

#--------EOF---------

MACRO ND3D2
  CLASS CORE ;
  FOREIGN ND3D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.544100 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 3.265 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 3.055 2.230 3.215 4.070 ;
        RECT 4.975 3.190 5.135 4.070 ;
        RECT 4.015 3.030 5.135 3.190 ;
        RECT 4.015 2.230 4.175 3.030 ;
        RECT 3.055 2.070 4.175 2.230 ;
        RECT 3.055 1.150 3.215 2.070 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.486200 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 2.505 2.085 3.680 2.215 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.590 2.720 2.000 ;
        RECT 3.550 1.590 3.680 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.486200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 1.590 1.760 4.000 ;
        RECT 4.510 1.590 4.640 4.000 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 3.945 0.475 4.245 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 1.630 0.345 4.640 0.475 ;
        RECT 3.945 0.260 4.245 0.345 ;
      LAYER Metal1 ;
        RECT 4.015 0.490 4.175 1.150 ;
        RECT 3.965 0.330 4.225 0.490 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.486200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 1.590 0.800 4.000 ;
        RECT 5.470 2.300 5.600 4.000 ;
        RECT 5.385 2.000 5.685 2.300 ;
        RECT 5.470 1.590 5.600 2.000 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 1.065 0.475 1.365 0.560 ;
        RECT 0.670 0.345 1.365 0.475 ;
        RECT 1.065 0.260 1.365 0.345 ;
      LAYER Metal1 ;
        RECT 5.405 2.070 5.665 2.230 ;
        RECT 5.455 1.570 5.615 2.070 ;
        RECT 3.535 1.410 5.615 1.570 ;
        RECT 3.535 0.490 3.695 1.410 ;
        RECT 1.085 0.330 3.695 0.490 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
END ND3D2

#--------EOF---------

MACRO ND3D4
  CLASS CORE ;
  FOREIGN ND3D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.947100 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 10.945 4.790 ;
        RECT 4.975 1.570 5.135 4.630 ;
        RECT 3.005 1.410 9.025 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.975000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 3.550 2.215 3.680 4.045 ;
        RECT 4.510 2.215 4.640 4.045 ;
        RECT 6.430 2.215 6.560 4.045 ;
        RECT 7.390 2.215 7.520 4.045 ;
        RECT 8.265 2.215 8.565 2.300 ;
        RECT 2.590 2.085 9.440 2.215 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 8.265 2.000 8.565 2.085 ;
        RECT 8.350 1.640 8.480 2.000 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
      LAYER Metal1 ;
        RECT 8.335 2.230 8.495 2.710 ;
        RECT 8.285 2.070 8.545 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.975000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 1.630 3.175 1.760 4.045 ;
        RECT 2.590 3.175 2.720 4.045 ;
        RECT 1.630 3.045 2.720 3.175 ;
        RECT 8.350 3.175 8.480 4.045 ;
        RECT 10.270 3.175 10.400 4.045 ;
        RECT 8.350 3.045 10.400 3.175 ;
        RECT 1.630 1.640 1.760 3.045 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 7.390 1.640 7.520 1.820 ;
        RECT 10.270 1.640 10.400 3.045 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 7.390 0.560 7.520 0.920 ;
        RECT 7.305 0.475 7.605 0.560 ;
        RECT 10.270 0.475 10.400 0.920 ;
        RECT 1.630 0.345 10.400 0.475 ;
        RECT 7.305 0.260 7.605 0.345 ;
      LAYER Metal1 ;
        RECT 7.375 0.490 7.535 1.150 ;
        RECT 7.325 0.330 7.585 0.490 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150150 ;
    PORT
      LAYER GatPoly ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 11.230 3.260 11.360 4.045 ;
        RECT 11.145 2.960 11.445 3.260 ;
      LAYER Metal1 ;
        RECT 11.215 3.190 11.375 4.230 ;
        RECT 11.165 3.030 11.425 3.190 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 11.695 5.130 11.855 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 0.670 3.865 0.800 4.045 ;
        RECT 5.470 3.865 5.600 4.045 ;
        RECT 9.310 3.865 9.440 4.045 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 5.470 1.640 5.600 1.820 ;
        RECT 6.430 1.640 6.560 1.820 ;
        RECT 11.230 1.640 11.360 1.820 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
  END
END ND3D4

#--------EOF---------

MACRO NR2D0
  CLASS CORE ;
  FOREIGN NR2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.637800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 4.970 2.305 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
    END
  END vdd
END NR2D0

#--------EOF---------

MACRO NR2D1
  CLASS CORE ;
  FOREIGN NR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.275600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 4.070 2.305 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
    END
  END vdd
END NR2D1

#--------EOF---------

MACRO NR2D2
  CLASS CORE ;
  FOREIGN NR2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.191200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 4.070 2.305 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 2.095 3.190 2.255 4.070 ;
        RECT 2.095 3.030 3.215 3.190 ;
        RECT 3.055 1.570 3.215 3.030 ;
        RECT 1.085 1.410 1.345 1.570 ;
        RECT 3.005 1.410 3.265 1.570 ;
    END
  END zn
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 0.585 2.085 3.680 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 3.260 1.760 4.000 ;
        RECT 1.545 3.175 1.845 3.260 ;
        RECT 2.590 3.175 2.720 4.000 ;
        RECT 1.545 3.045 2.720 3.175 ;
        RECT 1.545 2.960 1.845 3.045 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 2.590 1.640 2.720 1.820 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 1.545 0.475 1.845 0.560 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 1.545 0.345 2.720 0.475 ;
        RECT 1.545 0.260 1.845 0.345 ;
      LAYER Metal1 ;
        RECT 1.565 3.030 1.825 3.190 ;
        RECT 1.615 0.490 1.775 3.030 ;
        RECT 1.565 0.330 1.825 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
END NR2D2

#--------EOF---------

MACRO NR2D4
  CLASS CORE ;
  FOREIGN NR2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.382400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 4.070 6.145 4.230 ;
        RECT 0.655 1.570 0.815 4.070 ;
        RECT 2.575 2.710 2.735 4.070 ;
        RECT 2.575 2.550 4.655 2.710 ;
        RECT 4.495 1.570 4.655 2.550 ;
        RECT 0.655 1.410 1.345 1.570 ;
        RECT 3.005 1.410 7.105 1.570 ;
    END
  END zn
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 4.640 5.775 ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 4.510 5.200 4.640 5.645 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.670 2.695 0.800 4.000 ;
        RECT 3.550 3.260 3.680 4.000 ;
        RECT 4.510 3.820 4.640 4.000 ;
        RECT 7.390 3.260 7.520 4.000 ;
        RECT 3.465 2.960 3.765 3.260 ;
        RECT 7.305 2.960 7.605 3.260 ;
        RECT 3.550 2.695 3.680 2.960 ;
        RECT 0.670 2.565 3.680 2.695 ;
        RECT 0.670 1.640 0.800 2.565 ;
        RECT 3.550 1.640 3.680 1.820 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 7.390 1.640 7.520 2.960 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 7.390 0.475 7.520 0.920 ;
        RECT 3.550 0.345 7.520 0.475 ;
      LAYER Metal1 ;
        RECT 3.485 3.030 7.585 3.190 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 3.260 1.760 4.000 ;
        RECT 1.545 3.175 1.845 3.260 ;
        RECT 2.590 3.175 2.720 4.000 ;
        RECT 1.545 3.045 2.720 3.175 ;
        RECT 1.545 2.960 1.845 3.045 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 1.545 2.085 6.560 2.215 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 3.030 1.825 3.190 ;
        RECT 1.615 2.230 1.775 3.030 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
END NR2D4

#--------EOF---------

MACRO NR3D0
  CLASS CORE ;
  FOREIGN NR3D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.180200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.135 1.410 3.215 1.570 ;
        RECT 1.135 1.150 1.295 1.410 ;
        RECT 3.055 1.150 3.215 1.410 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
    END
  END vdd
END NR3D0

#--------EOF---------

MACRO NR3D1
  CLASS CORE ;
  FOREIGN NR3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.000400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.575 4.070 3.265 4.230 ;
        RECT 2.575 1.570 2.735 4.070 ;
        RECT 1.085 1.410 3.265 1.570 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 5.470 3.260 5.600 4.000 ;
        RECT 2.025 3.175 2.325 3.260 ;
        RECT 0.670 3.045 2.325 3.175 ;
        RECT 0.670 1.640 0.800 3.045 ;
        RECT 2.025 2.960 2.325 3.045 ;
        RECT 5.385 2.960 5.685 3.260 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 2.095 4.630 5.615 4.790 ;
        RECT 2.095 3.190 2.255 4.630 ;
        RECT 5.455 3.190 5.615 4.630 ;
        RECT 2.045 3.030 2.305 3.190 ;
        RECT 5.405 3.030 5.665 3.190 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 3.820 1.760 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 1.545 2.695 1.845 2.780 ;
        RECT 3.465 2.695 3.765 2.780 ;
        RECT 1.545 2.565 3.765 2.695 ;
        RECT 1.545 2.480 1.845 2.565 ;
        RECT 3.465 2.480 3.765 2.565 ;
        RECT 1.630 1.640 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 1.615 2.710 1.775 5.630 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 4.495 2.710 4.655 3.030 ;
        RECT 1.565 2.550 1.825 2.710 ;
        RECT 3.485 2.550 4.655 2.710 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.590 3.175 2.720 4.000 ;
        RECT 3.550 3.175 3.680 4.000 ;
        RECT 2.590 3.045 4.160 3.175 ;
        RECT 2.985 2.215 3.285 2.300 ;
        RECT 4.030 2.215 4.160 3.045 ;
        RECT 2.590 2.085 4.160 2.215 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 2.985 2.000 3.285 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 3.055 2.230 3.215 2.710 ;
        RECT 3.005 2.070 3.265 2.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
END NR3D1

#--------EOF---------

MACRO NR3D2
  CLASS CORE ;
  FOREIGN NR3D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.260 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.784800 ;
    PORT
      LAYER Metal1 ;
        RECT 9.725 4.070 11.905 4.230 ;
        RECT 9.775 1.570 9.935 4.070 ;
        RECT 3.005 1.410 9.985 1.570 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.811200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 0.670 3.045 1.760 3.175 ;
        RECT 1.630 2.215 1.760 3.045 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 1.630 2.085 3.680 2.215 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.811200 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 5.470 2.215 5.600 3.045 ;
        RECT 6.430 2.300 6.560 4.000 ;
        RECT 6.345 2.215 6.645 2.300 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 5.470 2.085 7.520 2.215 ;
        RECT 6.345 2.000 6.645 2.085 ;
        RECT 6.430 1.640 6.560 2.000 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 6.415 2.230 6.575 2.710 ;
        RECT 6.365 2.070 6.625 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.811200 ;
    PORT
      LAYER GatPoly ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 9.310 2.300 9.440 4.000 ;
        RECT 10.270 3.175 10.400 4.000 ;
        RECT 11.230 3.175 11.360 4.000 ;
        RECT 12.190 3.175 12.320 4.000 ;
        RECT 10.270 3.045 12.320 3.175 ;
        RECT 9.225 2.215 9.525 2.300 ;
        RECT 10.270 2.215 10.400 3.045 ;
        RECT 9.225 2.085 10.400 2.215 ;
        RECT 9.225 2.000 9.525 2.085 ;
        RECT 9.310 1.640 9.440 2.000 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
      LAYER Metal1 ;
        RECT 9.295 2.230 9.455 2.710 ;
        RECT 9.245 2.070 9.505 2.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 4.925 4.630 12.865 4.790 ;
        RECT 0.125 4.070 8.065 4.230 ;
  END
END NR3D2

#--------EOF---------

MACRO NR3D4
  CLASS CORE ;
  FOREIGN NR3D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.820 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.569600 ;
    PORT
      LAYER Metal1 ;
        RECT 17.405 4.070 17.665 4.230 ;
        RECT 19.325 4.070 23.425 4.230 ;
        RECT 17.455 1.570 17.615 4.070 ;
        RECT 19.375 1.570 19.535 4.070 ;
        RECT 4.925 1.410 19.585 1.570 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.622400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 0.670 3.045 1.760 3.175 ;
        RECT 1.630 2.215 1.760 3.045 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 1.630 2.085 7.520 2.215 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.622400 ;
    PORT
      LAYER GatPoly ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 8.350 3.175 8.480 4.000 ;
        RECT 9.310 3.175 9.440 4.000 ;
        RECT 8.350 3.045 9.440 3.175 ;
        RECT 9.310 2.215 9.440 3.045 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.300 12.320 4.000 ;
        RECT 12.105 2.215 12.405 2.300 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 14.110 2.215 14.240 4.000 ;
        RECT 15.070 2.215 15.200 4.000 ;
        RECT 9.310 2.085 15.200 2.215 ;
        RECT 12.105 2.000 12.405 2.085 ;
        RECT 12.190 1.640 12.320 2.000 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 14.110 1.640 14.240 2.085 ;
        RECT 15.070 1.640 15.200 2.085 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
      LAYER Metal1 ;
        RECT 12.175 2.230 12.335 2.710 ;
        RECT 12.125 2.070 12.385 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.622400 ;
    PORT
      LAYER GatPoly ;
        RECT 16.990 5.200 17.120 5.380 ;
        RECT 17.950 5.200 18.080 5.380 ;
        RECT 18.910 5.200 19.040 5.380 ;
        RECT 19.870 5.200 20.000 5.380 ;
        RECT 20.830 5.200 20.960 5.380 ;
        RECT 21.790 5.200 21.920 5.380 ;
        RECT 22.750 5.200 22.880 5.380 ;
        RECT 23.710 5.200 23.840 5.380 ;
        RECT 16.990 2.300 17.120 4.000 ;
        RECT 16.905 2.215 17.205 2.300 ;
        RECT 17.950 2.215 18.080 4.000 ;
        RECT 18.910 2.215 19.040 4.000 ;
        RECT 19.870 3.175 20.000 4.000 ;
        RECT 20.830 3.175 20.960 4.000 ;
        RECT 21.790 3.175 21.920 4.000 ;
        RECT 22.750 3.175 22.880 4.000 ;
        RECT 23.710 3.175 23.840 4.000 ;
        RECT 19.870 3.045 23.840 3.175 ;
        RECT 19.870 2.215 20.000 3.045 ;
        RECT 16.905 2.085 20.000 2.215 ;
        RECT 16.905 2.000 17.205 2.085 ;
        RECT 16.990 1.640 17.120 2.000 ;
        RECT 17.950 1.640 18.080 2.085 ;
        RECT 18.910 1.640 19.040 2.085 ;
        RECT 19.870 1.640 20.000 2.085 ;
        RECT 16.990 0.740 17.120 0.920 ;
        RECT 17.950 0.740 18.080 0.920 ;
        RECT 18.910 0.740 19.040 0.920 ;
        RECT 19.870 0.740 20.000 0.920 ;
      LAYER Metal1 ;
        RECT 16.975 2.230 17.135 2.710 ;
        RECT 16.925 2.070 17.185 2.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 15.485 0.990 15.745 1.150 ;
        RECT 16.445 0.990 16.705 1.150 ;
        RECT 18.365 0.990 18.625 1.150 ;
        RECT 20.285 0.990 20.545 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 15.535 0.150 15.695 0.990 ;
        RECT 16.495 0.150 16.655 0.990 ;
        RECT 18.415 0.150 18.575 0.990 ;
        RECT 20.335 0.150 20.495 0.990 ;
        RECT 0.000 -0.150 24.820 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 24.820 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 8.765 4.630 24.385 4.790 ;
        RECT 0.125 4.070 15.745 4.230 ;
  END
END NR3D4

#--------EOF---------

MACRO OA21D0
  CLASS CORE ;
  FOREIGN OA21D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 2.590 2.215 2.720 4.600 ;
        RECT 2.025 2.085 2.720 2.215 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 2.590 1.280 2.720 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.095 2.230 2.255 2.710 ;
        RECT 2.045 2.070 2.305 2.230 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 1.150 4.175 4.970 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.600 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.280 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.970 2.735 5.130 ;
        RECT 2.575 2.230 2.735 4.970 ;
        RECT 2.575 2.070 3.745 2.230 ;
        RECT 0.655 1.410 2.255 1.570 ;
        RECT 0.655 1.150 0.815 1.410 ;
        RECT 2.095 1.150 2.255 1.410 ;
        RECT 2.575 1.150 2.735 2.070 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 1.085 0.990 2.735 1.150 ;
  END
END OA21D0

#--------EOF---------

MACRO OA21D1
  CLASS CORE ;
  FOREIGN OA21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 3.965 1.410 4.225 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 3.485 2.070 3.745 2.230 ;
        RECT 3.535 1.570 3.695 2.070 ;
        RECT 1.085 1.410 3.695 1.570 ;
        RECT 0.125 0.990 2.305 1.150 ;
  END
END OA21D1

#--------EOF---------

MACRO OA21D2
  CLASS CORE ;
  FOREIGN OA21D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.000 4.725 2.300 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 0.670 2.085 1.845 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 1.615 1.570 1.775 2.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.615 1.410 4.225 1.570 ;
        RECT 3.005 0.990 5.185 1.150 ;
  END
END OA21D2

#--------EOF---------

MACRO OA21D4
  CLASS CORE ;
  FOREIGN OA21D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.540 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 0.670 3.045 1.760 3.175 ;
        RECT 1.630 2.215 1.760 3.045 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 4.510 2.215 4.640 3.045 ;
        RECT 1.630 2.085 4.640 2.215 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 4.425 5.560 4.725 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 4.510 5.200 4.640 5.560 ;
        RECT 1.630 3.820 1.760 4.000 ;
        RECT 4.510 3.820 4.640 4.000 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.475 4.725 0.560 ;
        RECT 1.630 0.345 4.725 0.475 ;
        RECT 4.425 0.260 4.725 0.345 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 4.445 5.630 4.705 5.790 ;
        RECT 1.615 4.790 1.775 5.630 ;
        RECT 4.495 4.790 4.655 5.630 ;
        RECT 1.615 4.630 4.655 4.790 ;
        RECT 4.495 0.490 4.655 4.630 ;
        RECT 4.445 0.330 4.705 0.490 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 3.260 3.680 4.000 ;
        RECT 3.465 2.960 3.765 3.260 ;
      LAYER Metal1 ;
        RECT 3.055 3.030 3.745 3.190 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 6.895 1.570 7.055 4.070 ;
        RECT 8.815 1.570 8.975 4.070 ;
        RECT 6.845 1.410 9.025 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 0.000 -0.150 10.540 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 10.540 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 2.590 3.820 2.720 4.000 ;
        RECT 6.430 3.820 6.560 4.000 ;
        RECT 7.390 3.820 7.520 4.000 ;
        RECT 8.350 3.820 8.480 4.000 ;
        RECT 9.310 3.820 9.440 4.000 ;
        RECT 0.670 1.640 0.800 1.820 ;
        RECT 5.470 1.640 5.600 1.820 ;
        RECT 6.430 1.640 6.560 1.820 ;
        RECT 7.390 1.640 7.520 1.820 ;
        RECT 8.350 1.640 8.480 1.820 ;
        RECT 9.310 1.640 9.440 1.820 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.070 4.225 4.230 ;
        RECT 4.015 1.150 4.175 4.070 ;
        RECT 2.045 0.990 4.225 1.150 ;
  END
END OA21D4

#--------EOF---------

MACRO OAI21D0
  CLASS CORE ;
  FOREIGN OAI21D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.796800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 1.135 4.630 2.255 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 1.615 0.990 2.305 1.150 ;
        RECT 1.615 0.490 1.775 0.990 ;
        RECT 0.655 0.330 1.775 0.490 ;
  END
END OAI21D0

#--------EOF---------

MACRO OAI21D1
  CLASS CORE ;
  FOREIGN OAI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 2.095 3.190 2.255 4.070 ;
        RECT 1.135 3.030 2.255 3.190 ;
        RECT 1.135 1.570 1.295 3.030 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 2.305 1.150 ;
  END
END OAI21D1

#--------EOF---------

MACRO OAI21D2
  CLASS CORE ;
  FOREIGN OAI21D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.070 4.225 4.230 ;
        RECT 4.015 1.150 4.175 4.070 ;
        RECT 2.045 0.990 4.225 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 1.630 3.045 2.720 3.175 ;
        RECT 2.590 2.300 2.720 3.045 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 4.510 2.215 4.640 4.000 ;
        RECT 2.505 2.085 4.640 2.215 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 4.510 1.640 4.640 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 0.670 2.695 0.800 4.000 ;
        RECT 5.470 3.260 5.600 4.000 ;
        RECT 5.385 2.960 5.685 3.260 ;
        RECT 0.670 2.565 1.760 2.695 ;
        RECT 1.630 1.640 1.760 2.565 ;
        RECT 3.550 1.640 3.680 1.820 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 3.465 0.475 3.765 0.560 ;
        RECT 1.630 0.345 3.765 0.475 ;
        RECT 3.465 0.260 3.765 0.345 ;
      LAYER Metal1 ;
        RECT 4.495 3.030 5.665 3.190 ;
        RECT 4.495 0.490 4.655 3.030 ;
        RECT 3.485 0.330 4.655 0.490 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 2.505 5.560 2.805 5.860 ;
        RECT 2.590 5.200 2.720 5.560 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.590 3.820 2.720 4.000 ;
        RECT 3.550 3.260 3.680 4.000 ;
        RECT 3.465 2.960 3.765 3.260 ;
        RECT 5.865 2.960 6.165 3.260 ;
        RECT 5.950 2.695 6.080 2.960 ;
        RECT 5.470 2.565 6.080 2.695 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 5.470 1.640 5.600 2.565 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 5.630 2.785 5.790 ;
        RECT 2.575 4.790 2.735 5.630 ;
        RECT 1.615 4.630 6.095 4.790 ;
        RECT 1.615 3.190 1.775 4.630 ;
        RECT 5.935 3.190 6.095 4.630 ;
        RECT 1.615 3.030 3.745 3.190 ;
        RECT 5.885 3.030 6.145 3.190 ;
        RECT 1.615 2.230 1.775 3.030 ;
        RECT 0.605 2.070 1.775 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
END OAI21D2

#--------EOF---------

MACRO OAI21D4
  CLASS CORE ;
  FOREIGN OAI21D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.260 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.176000 ;
    PORT
      LAYER GatPoly ;
        RECT 8.265 2.480 8.565 2.780 ;
        RECT 8.350 1.640 8.480 2.480 ;
        RECT 8.265 1.340 8.565 1.640 ;
      LAYER Metal1 ;
        RECT 1.085 4.070 3.265 4.230 ;
        RECT 9.725 4.070 11.905 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 9.775 3.190 9.935 4.070 ;
        RECT 8.815 3.030 9.935 3.190 ;
        RECT 7.375 2.550 8.545 2.710 ;
        RECT 7.375 1.570 7.535 2.550 ;
        RECT 8.815 2.230 8.975 3.030 ;
        RECT 1.085 1.410 7.535 1.570 ;
        RECT 7.855 2.070 8.975 2.230 ;
        RECT 1.135 1.150 1.295 1.410 ;
        RECT 7.855 1.150 8.015 2.070 ;
        RECT 8.285 1.410 11.905 1.570 ;
        RECT 0.125 0.990 8.065 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 0.585 2.085 3.680 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 7.390 3.175 7.520 4.000 ;
        RECT 8.350 3.175 8.480 4.000 ;
        RECT 7.390 3.045 8.480 3.175 ;
        RECT 7.390 2.215 7.520 3.045 ;
        RECT 4.425 2.085 7.520 2.215 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.085 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 9.310 2.300 9.440 4.000 ;
        RECT 9.225 2.215 9.525 2.300 ;
        RECT 10.270 2.215 10.400 4.000 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 9.225 2.085 12.320 2.215 ;
        RECT 9.225 2.000 9.525 2.085 ;
        RECT 9.310 1.640 9.440 2.000 ;
        RECT 10.270 1.640 10.400 2.085 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
      LAYER Metal1 ;
        RECT 9.295 2.230 9.455 2.710 ;
        RECT 9.245 2.070 9.505 2.230 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 12.655 0.150 12.815 0.990 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 12.655 5.130 12.815 5.970 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 8.065 4.790 ;
  END
END OAI21D4

#--------EOF---------

MACRO OAI211D0
  CLASS CORE ;
  FOREIGN OAI211D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.600 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.280 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.600 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.280 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END c
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 4.015 4.790 4.175 4.970 ;
        RECT 1.135 4.630 4.175 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 1.615 0.990 2.305 1.150 ;
        RECT 1.615 0.490 1.775 0.990 ;
        RECT 0.655 0.330 1.775 0.490 ;
  END
END OAI211D0

#--------EOF---------

MACRO OAI211D1
  CLASS CORE ;
  FOREIGN OAI211D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.000 2.805 2.300 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END c
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.271600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.070 4.225 4.230 ;
        RECT 2.095 3.190 2.255 4.070 ;
        RECT 1.135 3.030 2.255 3.190 ;
        RECT 1.135 1.570 1.295 3.030 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 2.305 1.150 ;
  END
END OAI211D1

#--------EOF---------

MACRO OAI211D2
  CLASS CORE ;
  FOREIGN OAI211D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 4.425 2.085 7.520 2.215 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 7.390 1.640 7.520 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 6.430 3.260 6.560 4.000 ;
        RECT 6.345 3.175 6.645 3.260 ;
        RECT 5.470 3.045 6.645 3.175 ;
        RECT 6.345 2.960 6.645 3.045 ;
        RECT 5.470 1.640 5.600 1.820 ;
        RECT 6.430 1.640 6.560 1.820 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 6.430 0.560 6.560 0.920 ;
        RECT 6.345 0.475 6.645 0.560 ;
        RECT 5.470 0.345 6.645 0.475 ;
        RECT 6.345 0.260 6.645 0.345 ;
      LAYER Metal1 ;
        RECT 6.365 3.030 6.625 3.190 ;
        RECT 6.415 0.490 6.575 3.030 ;
        RECT 6.365 0.330 6.625 0.490 ;
    END
  END c
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.192000 ;
    PORT
      LAYER GatPoly ;
        RECT 5.865 2.695 6.165 2.780 ;
        RECT 6.825 2.695 7.125 2.780 ;
        RECT 5.865 2.565 7.125 2.695 ;
        RECT 5.865 2.480 6.165 2.565 ;
        RECT 6.825 2.480 7.125 2.565 ;
      LAYER Metal1 ;
        RECT 1.615 4.630 7.535 4.790 ;
        RECT 1.615 2.710 1.775 4.630 ;
        RECT 2.045 4.070 7.105 4.230 ;
        RECT 0.655 2.550 1.775 2.710 ;
        RECT 0.655 1.570 0.815 2.550 ;
        RECT 0.125 1.410 0.815 1.570 ;
        RECT 1.615 1.570 1.775 2.550 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 7.375 2.710 7.535 4.630 ;
        RECT 5.885 2.550 6.145 2.710 ;
        RECT 6.845 2.550 8.015 2.710 ;
        RECT 5.935 1.570 6.095 2.550 ;
        RECT 7.855 1.570 8.015 2.550 ;
        RECT 1.615 1.410 2.305 1.570 ;
        RECT 3.965 1.410 6.095 1.570 ;
        RECT 7.805 1.410 8.065 1.570 ;
        RECT 2.095 1.150 2.255 1.410 ;
        RECT 1.085 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.065 2.215 1.365 2.300 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 0.670 2.085 3.680 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.065 2.000 1.365 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 2.070 1.345 2.230 ;
        RECT 1.135 1.410 1.295 2.070 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499200 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 2.590 3.260 2.720 4.000 ;
        RECT 2.505 3.175 2.805 3.260 ;
        RECT 1.630 3.045 2.805 3.175 ;
        RECT 2.505 2.960 2.805 3.045 ;
        RECT 1.630 1.640 1.760 1.820 ;
        RECT 2.590 1.640 2.720 1.820 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 3.465 0.475 3.765 0.560 ;
        RECT 1.630 0.345 3.765 0.475 ;
        RECT 3.465 0.260 3.765 0.345 ;
      LAYER Metal1 ;
        RECT 2.525 3.030 3.695 3.190 ;
        RECT 3.535 0.490 3.695 3.030 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
END OAI211D2

#--------EOF---------

MACRO OAI211D4
  CLASS CORE ;
  FOREIGN OAI211D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.000 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.582399 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 15.745 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 0.125 1.410 8.065 1.570 ;
    END
  END zn
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 0.670 2.085 3.680 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
#        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.560 2.070 1.84 2.710 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.645 8.480 5.775 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 6.430 5.200 6.560 5.645 ;
        RECT 7.390 5.200 7.520 5.645 ;
        RECT 8.350 5.200 8.480 5.645 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 4.510 1.640 4.640 3.045 ;
        RECT 5.470 1.640 5.600 3.045 ;
        RECT 6.430 1.640 6.560 4.000 ;
        RECT 7.390 2.300 7.520 4.000 ;
        RECT 8.350 3.820 8.480 4.000 ;
        RECT 7.305 2.000 7.605 2.300 ;
        RECT 7.390 1.640 7.520 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
#        RECT 7.375 2.230 7.535 2.710 ;
        RECT 7.320 2.070 7.600 2.710 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 9.310 2.695 9.440 4.000 ;
        RECT 10.270 2.695 10.400 4.000 ;
        RECT 11.230 2.780 11.360 4.000 ;
        RECT 11.145 2.695 11.445 2.780 ;
        RECT 12.190 2.695 12.320 4.000 ;
        RECT 9.310 2.565 12.320 2.695 ;
        RECT 9.310 1.640 9.440 2.565 ;
        RECT 10.270 1.640 10.400 2.565 ;
        RECT 11.145 2.480 11.445 2.565 ;
        RECT 11.230 1.640 11.360 2.480 ;
        RECT 12.190 1.640 12.320 2.565 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
      LAYER Metal1 ;
#        RECT 11.215 2.710 11.375 3.190 ;
        RECT 11.160 2.550 11.440 3.190 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.998400 ;
    PORT
      LAYER GatPoly ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 16.030 5.200 16.160 5.380 ;
        RECT 13.150 3.260 13.280 4.000 ;
        RECT 13.065 3.175 13.365 3.260 ;
        RECT 14.110 3.175 14.240 4.000 ;
        RECT 15.070 3.175 15.200 4.000 ;
        RECT 16.030 3.175 16.160 4.000 ;
        RECT 13.065 3.045 16.160 3.175 ;
        RECT 13.065 2.960 13.365 3.045 ;
        RECT 13.150 1.640 13.280 2.960 ;
        RECT 14.110 1.640 14.240 3.045 ;
        RECT 15.070 1.640 15.200 3.045 ;
        RECT 16.030 1.640 16.160 3.045 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
        RECT 16.030 0.740 16.160 0.920 ;
      LAYER Metal1 ;
        RECT 13.080 2.550 13.36 3.190 ;
#        RECT 13.135 2.550 13.295 3.030 ;
    END
  END c
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 15.485 0.990 15.745 1.150 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 15.535 0.150 15.695 0.990 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 17.000 6.270 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 12.655 5.130 12.815 5.970 ;
        RECT 14.575 5.130 14.735 5.970 ;
        RECT 16.495 5.130 16.655 5.970 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 14.525 4.970 14.785 5.130 ;
        RECT 16.445 4.970 16.705 5.130 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 8.065 4.790 ;
        RECT 8.765 1.410 16.705 1.570 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 11.905 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OAI211D4

#--------EOF---------

MACRO OR2D0
  CLASS CORE ;
  FOREIGN OR2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 1.150 3.215 4.970 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.780 1.760 4.600 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 1.280 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.710 1.775 3.190 ;
        RECT 1.565 2.550 1.825 2.710 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 2.590 2.215 2.720 4.600 ;
        RECT 2.025 2.085 2.720 2.215 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 2.590 1.280 2.720 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 0.175 4.630 1.295 4.790 ;
        RECT 1.135 2.230 1.295 4.630 ;
        RECT 1.135 2.070 2.305 2.230 ;
        RECT 1.135 1.150 1.295 2.070 ;
        RECT 1.085 0.990 1.345 1.150 ;
  END
END OR2D0

#--------EOF---------

MACRO OR2D1
  CLASS CORE ;
  FOREIGN OR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.048075 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.241150 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.575 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.241150 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.780 1.760 4.000 ;
        RECT 1.545 2.480 1.845 2.780 ;
        RECT 1.630 1.575 1.760 2.480 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.710 1.775 3.190 ;
        RECT 1.565 2.550 1.825 2.710 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 2.025 2.085 2.720 2.215 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 2.590 1.575 2.720 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 3.190 0.335 4.070 ;
        RECT 0.175 3.030 1.295 3.190 ;
        RECT 1.135 2.230 1.295 3.030 ;
        RECT 1.135 2.070 2.305 2.230 ;
        RECT 1.135 1.150 1.295 2.070 ;
        RECT 1.085 0.990 1.345 1.150 ;
  END
END OR2D1

#--------EOF---------

MACRO OR2D2
  CLASS CORE ;
  FOREIGN OR2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 1.085 1.410 1.345 1.570 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202800 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 3.550 1.280 3.680 2.000 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.230 3.695 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202800 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.780 2.720 4.000 ;
        RECT 2.505 2.480 2.805 2.780 ;
        RECT 2.590 1.280 2.720 2.480 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.710 2.735 3.190 ;
        RECT 2.525 2.550 2.785 2.710 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 0.670 2.085 2.325 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 4.015 3.190 4.175 4.070 ;
        RECT 3.055 3.030 4.175 3.190 ;
        RECT 3.055 2.230 3.215 3.030 ;
        RECT 2.045 2.070 3.215 2.230 ;
        RECT 3.055 1.150 3.215 2.070 ;
        RECT 3.005 0.990 3.265 1.150 ;
  END
END OR2D2

#--------EOF---------

MACRO OR2D4
  CLASS CORE ;
  FOREIGN OR2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.070 1.345 4.230 ;
        RECT 3.005 4.070 3.265 4.230 ;
        RECT 1.135 1.570 1.295 4.070 ;
        RECT 3.055 1.570 3.215 4.070 ;
        RECT 1.085 1.410 3.265 1.570 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405600 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 5.865 3.175 6.165 3.260 ;
        RECT 6.430 3.175 6.560 4.000 ;
        RECT 5.470 3.045 6.560 3.175 ;
        RECT 5.470 1.555 5.600 3.045 ;
        RECT 5.865 2.960 6.165 3.045 ;
        RECT 5.470 1.425 6.560 1.555 ;
        RECT 5.470 1.280 5.600 1.425 ;
        RECT 6.430 1.280 6.560 1.425 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 5.885 3.030 6.145 3.190 ;
        RECT 5.935 2.550 6.095 3.030 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 4.510 1.555 4.640 4.000 ;
        RECT 7.390 2.300 7.520 4.000 ;
        RECT 4.905 2.000 5.205 2.300 ;
        RECT 7.305 2.000 7.605 2.300 ;
        RECT 4.990 1.555 5.120 2.000 ;
        RECT 4.510 1.425 5.120 1.555 ;
        RECT 4.510 1.280 4.640 1.425 ;
        RECT 7.390 1.280 7.520 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
      LAYER Metal1 ;
        RECT 4.925 2.070 7.585 2.230 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 7.855 0.150 8.015 0.990 ;
        RECT 0.000 -0.150 8.500 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 8.500 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 2.095 5.130 2.255 5.970 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 7.855 5.130 8.015 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.215 2.720 4.000 ;
        RECT 3.550 2.215 3.680 4.000 ;
        RECT 3.945 2.215 4.245 2.300 ;
        RECT 0.670 2.085 4.245 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.590 1.640 2.720 2.085 ;
        RECT 3.550 1.640 3.680 2.085 ;
        RECT 3.945 2.000 4.245 2.085 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 5.455 4.070 6.145 4.230 ;
        RECT 5.455 2.710 5.615 4.070 ;
        RECT 4.495 2.550 5.615 2.710 ;
        RECT 4.495 2.230 4.655 2.550 ;
        RECT 3.965 2.070 4.655 2.230 ;
        RECT 4.495 1.570 4.655 2.070 ;
        RECT 4.495 1.410 7.055 1.570 ;
        RECT 4.975 1.150 5.135 1.410 ;
        RECT 6.895 1.150 7.055 1.410 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
  END
END OR2D4

#--------EOF---------

MACRO TAPCELL
  CLASS CORE ;
  FOREIGN TAPCELL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.380 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.590 0.920 0.850 1.080 ;
        RECT 1.070 0.920 1.330 1.080 ;
        RECT 1.550 0.920 1.810 1.080 ;
        RECT 0.640 0.150 0.800 0.920 ;
        RECT 1.120 0.150 1.280 0.920 ;
        RECT 1.600 0.150 1.760 0.920 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.380 6.270 ;
        RECT 0.640 5.200 0.800 5.970 ;
        RECT 1.120 5.200 1.280 5.970 ;
        RECT 1.600 5.200 1.760 5.970 ;
        RECT 0.590 5.040 0.850 5.200 ;
        RECT 1.070 5.040 1.330 5.200 ;
        RECT 1.550 5.040 1.810 5.200 ;
    END
  END vdd
END TAPCELL

#--------EOF---------

MACRO TIEH
  CLASS CORE ;
  FOREIGN TIEH ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 4.070 0.335 5.130 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 1.640 0.800 4.000 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH

#--------EOF---------

MACRO TIEL
  CLASS CORE ;
  FOREIGN TIEL ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.990 0.335 2.230 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.105 3.175 0.405 3.260 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 0.105 3.045 0.800 3.175 ;
        RECT 0.105 2.960 0.405 3.045 ;
        RECT 0.670 1.640 0.800 3.045 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 3.190 0.335 4.070 ;
        RECT 0.125 3.030 0.385 3.190 ;
  END
END TIEL

#--------EOF---------

MACRO XNR2D0
  CLASS CORE ;
  FOREIGN XNR2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.170300 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 5.600 5.775 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 3.550 4.615 3.680 4.795 ;
        RECT 2.590 1.170 2.720 1.350 ;
        RECT 5.470 1.170 5.600 4.795 ;
        RECT 2.590 0.560 2.720 0.920 ;
        RECT 2.505 0.475 2.805 0.560 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 2.505 0.345 5.600 0.475 ;
        RECT 2.505 0.260 2.805 0.345 ;
      LAYER Metal1 ;
        RECT 2.575 0.490 2.735 1.150 ;
        RECT 2.525 0.330 2.785 0.490 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.300 1.760 4.600 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.280 1.760 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.230 1.775 2.710 ;
        RECT 1.565 2.070 1.825 2.230 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 0.670 3.260 0.800 4.600 ;
        RECT 2.025 4.000 2.325 4.300 ;
        RECT 2.590 4.215 2.720 4.795 ;
        RECT 3.945 4.215 4.245 4.300 ;
        RECT 2.590 4.085 4.245 4.215 ;
        RECT 3.945 4.000 4.245 4.085 ;
        RECT 0.585 2.960 0.885 3.260 ;
        RECT 2.110 3.175 2.240 4.000 ;
        RECT 4.510 3.175 4.640 4.795 ;
        RECT 2.110 3.045 5.120 3.175 ;
        RECT 0.670 1.280 0.800 2.960 ;
        RECT 2.110 2.300 2.240 3.045 ;
        RECT 2.025 2.000 2.325 2.300 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 3.550 2.085 4.725 2.215 ;
        RECT 3.550 1.170 3.680 2.085 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.990 1.555 5.120 3.045 ;
        RECT 4.510 1.425 5.120 1.555 ;
        RECT 4.510 1.170 4.640 1.425 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 5.455 4.970 6.145 5.130 ;
        RECT 2.095 4.230 2.255 4.970 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.055 3.190 3.215 4.970 ;
        RECT 0.605 3.030 3.215 3.190 ;
        RECT 2.045 2.070 2.305 2.230 ;
        RECT 2.095 1.150 2.255 2.070 ;
        RECT 3.055 1.150 3.215 3.030 ;
        RECT 3.535 1.150 3.695 4.970 ;
        RECT 5.455 4.230 5.615 4.970 ;
        RECT 3.965 4.070 6.095 4.230 ;
        RECT 5.455 2.230 5.615 4.070 ;
        RECT 5.935 2.230 6.095 4.070 ;
        RECT 4.445 2.070 6.095 2.230 ;
        RECT 5.935 1.150 6.095 2.070 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.535 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
  END
END XNR2D0

#--------EOF---------

MACRO XNR2D1
  CLASS CORE ;
  FOREIGN XNR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.175 1.760 4.000 ;
        RECT 2.025 3.175 2.325 3.260 ;
        RECT 1.630 3.045 2.325 3.175 ;
        RECT 2.025 2.960 2.325 3.045 ;
        RECT 2.025 2.215 2.325 2.300 ;
        RECT 1.630 2.085 2.325 2.215 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.025 2.000 2.325 2.085 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 3.030 2.305 3.190 ;
        RECT 2.095 2.230 2.255 3.030 ;
        RECT 2.045 2.070 2.305 2.230 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 5.885 1.410 6.145 1.570 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 4.300 0.800 4.600 ;
        RECT 0.585 4.000 0.885 4.300 ;
        RECT 2.985 4.215 3.285 4.300 ;
        RECT 3.550 4.215 3.680 4.600 ;
        RECT 2.985 4.085 3.680 4.215 ;
        RECT 2.985 4.000 3.285 4.085 ;
        RECT 3.070 1.555 3.200 4.000 ;
        RECT 0.670 1.280 0.800 1.460 ;
        RECT 2.590 1.425 3.200 1.555 ;
        RECT 2.590 1.280 2.720 1.425 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 0.670 0.345 2.720 0.475 ;
      LAYER Metal1 ;
        RECT 0.655 4.630 2.735 4.790 ;
        RECT 0.655 4.230 0.815 4.630 ;
        RECT 2.575 4.230 2.735 4.630 ;
        RECT 0.605 4.070 0.865 4.230 ;
        RECT 2.575 4.070 3.265 4.230 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.425 5.560 4.725 5.860 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.560 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 2.590 2.780 2.720 4.600 ;
        RECT 4.510 4.420 4.640 4.600 ;
        RECT 3.945 3.175 4.245 3.260 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 3.945 3.045 5.600 3.175 ;
        RECT 3.945 2.960 4.245 3.045 ;
        RECT 0.105 2.695 0.405 2.780 ;
        RECT 2.505 2.695 2.805 2.780 ;
        RECT 0.105 2.565 2.805 2.695 ;
        RECT 0.105 2.480 0.405 2.565 ;
        RECT 2.505 2.480 2.805 2.565 ;
        RECT 3.465 2.480 3.765 2.780 ;
        RECT 3.550 1.280 3.680 2.480 ;
        RECT 3.945 2.215 4.245 2.300 ;
        RECT 5.470 2.215 5.600 3.045 ;
        RECT 3.945 2.085 5.600 2.215 ;
        RECT 3.945 2.000 4.245 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 4.510 1.280 4.640 1.460 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 4.425 0.260 4.725 0.560 ;
      LAYER Metal1 ;
        RECT 2.575 5.630 4.705 5.790 ;
        RECT 2.575 5.130 2.735 5.630 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.735 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.965 4.970 4.655 5.130 ;
        RECT 0.175 2.710 0.335 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 3.055 4.630 4.175 4.790 ;
        RECT 1.615 4.070 2.305 4.230 ;
        RECT 0.125 2.550 0.385 2.710 ;
        RECT 0.175 1.150 0.335 2.550 ;
        RECT 1.615 1.570 1.775 4.070 ;
        RECT 4.015 3.190 4.175 4.630 ;
        RECT 3.965 3.030 4.225 3.190 ;
        RECT 2.525 2.550 3.745 2.710 ;
        RECT 3.535 2.070 4.225 2.230 ;
        RECT 1.615 1.410 2.305 1.570 ;
        RECT 3.535 1.150 3.695 2.070 ;
        RECT 4.495 1.150 4.655 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.735 1.150 ;
        RECT 3.005 0.990 3.695 1.150 ;
        RECT 3.965 0.990 4.655 1.150 ;
        RECT 2.575 0.490 2.735 0.990 ;
        RECT 2.575 0.330 4.705 0.490 ;
  END
END XNR2D1

#--------EOF---------

MACRO XNR2D2
  CLASS CORE ;
  FOREIGN XNR2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 0.670 3.175 0.800 4.600 ;
        RECT 2.590 3.175 2.720 4.600 ;
        RECT 0.670 3.045 2.720 3.175 ;
        RECT 0.670 1.280 0.800 3.045 ;
        RECT 3.550 1.280 3.680 1.460 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 3.465 0.475 3.765 0.560 ;
        RECT 0.670 0.345 3.765 0.475 ;
        RECT 3.465 0.260 3.765 0.345 ;
      LAYER Metal1 ;
        RECT 3.535 0.490 3.695 1.150 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 4.510 1.640 4.640 1.820 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.260 4.725 0.560 ;
      LAYER Metal1 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 4.495 0.490 4.655 3.030 ;
        RECT 4.445 0.330 4.705 0.490 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 5.885 1.410 6.145 1.570 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 3.820 1.760 4.000 ;
        RECT 1.065 2.695 1.365 2.780 ;
        RECT 3.550 2.695 3.680 4.600 ;
        RECT 1.065 2.565 3.680 2.695 ;
        RECT 5.470 3.175 5.600 4.000 ;
        RECT 6.430 3.175 6.560 4.000 ;
        RECT 5.470 3.045 6.560 3.175 ;
        RECT 5.470 2.695 5.600 3.045 ;
        RECT 5.470 2.565 6.560 2.695 ;
        RECT 1.065 2.480 1.365 2.565 ;
        RECT 1.545 2.000 1.845 2.300 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 2.590 1.280 2.720 2.565 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 5.470 2.215 5.600 2.565 ;
        RECT 3.465 2.085 5.600 2.215 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.430 1.640 6.560 2.565 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 2.575 5.630 3.695 5.790 ;
        RECT 1.615 5.130 1.775 5.630 ;
        RECT 2.575 5.130 2.735 5.630 ;
        RECT 3.535 5.130 3.695 5.630 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.615 4.970 2.735 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 0.175 4.630 1.295 4.790 ;
        RECT 1.135 2.710 1.295 4.630 ;
        RECT 1.085 2.550 1.345 2.710 ;
        RECT 1.135 2.230 1.295 2.550 ;
        RECT 1.615 2.230 1.775 4.970 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 0.175 2.070 1.295 2.230 ;
        RECT 1.565 2.070 1.825 2.230 ;
        RECT 0.175 1.150 0.335 2.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 3.055 2.230 3.215 4.970 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 3.055 2.070 3.745 2.230 ;
        RECT 2.045 1.410 2.305 1.570 ;
        RECT 3.055 1.150 3.215 2.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 3.965 1.410 4.225 1.570 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
  END
END XNR2D2

#--------EOF---------

MACRO XNR2D4
  CLASS CORE ;
  FOREIGN XNR2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.713700 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 4.510 3.175 4.640 4.000 ;
        RECT 4.510 3.045 5.600 3.175 ;
        RECT 5.470 2.300 5.600 3.045 ;
        RECT 5.385 2.215 5.685 2.300 ;
        RECT 7.390 2.215 7.520 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 5.385 2.085 9.440 2.215 ;
        RECT 5.385 2.000 5.685 2.085 ;
        RECT 5.470 1.505 5.600 2.000 ;
        RECT 6.430 1.505 6.560 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
      LAYER Metal1 ;
        RECT 5.455 2.230 5.615 2.710 ;
        RECT 5.405 2.070 5.665 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.748800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 0.670 2.085 2.805 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 10.685 4.070 10.945 4.230 ;
        RECT 12.605 4.070 12.865 4.230 ;
        RECT 10.735 1.570 10.895 4.070 ;
        RECT 12.655 1.570 12.815 4.070 ;
        RECT 10.685 1.410 12.865 1.570 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 11.695 5.130 11.855 5.970 ;
        RECT 13.615 5.130 13.775 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
        RECT 13.565 4.970 13.825 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 6.345 5.775 6.645 5.860 ;
        RECT 5.470 5.645 6.645 5.775 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 6.345 5.560 6.645 5.645 ;
        RECT 6.430 5.200 6.560 5.560 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 5.470 3.820 5.600 4.000 ;
        RECT 6.430 3.820 6.560 4.000 ;
        RECT 10.270 2.300 10.400 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 10.185 2.215 10.485 2.300 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 10.185 2.085 13.280 2.215 ;
        RECT 10.185 2.000 10.485 2.085 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 4.510 1.505 4.640 1.685 ;
        RECT 7.390 1.505 7.520 1.685 ;
        RECT 10.270 1.640 10.400 2.000 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 8.265 1.340 8.565 1.640 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 7.390 0.475 7.520 0.920 ;
        RECT 8.350 0.475 8.480 1.340 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 4.510 0.345 8.480 0.475 ;
      LAYER Metal1 ;
        RECT 6.365 5.630 6.625 5.790 ;
        RECT 6.415 5.130 6.575 5.630 ;
        RECT 6.415 4.970 8.495 5.130 ;
        RECT 4.495 4.630 8.065 4.790 ;
        RECT 4.495 4.230 4.655 4.630 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 3.965 4.070 4.655 4.230 ;
        RECT 4.925 4.070 5.185 4.230 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 6.845 4.070 7.105 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 3.485 2.070 3.745 2.230 ;
        RECT 3.535 1.570 3.695 2.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 0.125 1.410 3.695 1.570 ;
        RECT 3.965 1.410 4.225 1.570 ;
        RECT 3.535 1.150 3.695 1.410 ;
        RECT 4.975 1.150 5.135 4.070 ;
        RECT 5.935 1.150 6.095 4.070 ;
        RECT 6.895 1.150 7.055 4.070 ;
        RECT 7.375 1.570 7.535 4.630 ;
        RECT 8.335 4.230 8.495 4.970 ;
        RECT 8.335 4.070 9.025 4.230 ;
        RECT 8.335 1.570 8.495 4.070 ;
        RECT 9.295 2.070 10.465 2.230 ;
        RECT 7.375 1.410 8.015 1.570 ;
        RECT 8.285 1.410 9.025 1.570 ;
        RECT 7.855 1.150 8.015 1.410 ;
        RECT 9.295 1.150 9.455 2.070 ;
        RECT 3.535 0.990 6.145 1.150 ;
        RECT 6.415 0.990 9.455 1.150 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 6.415 0.490 6.575 0.990 ;
        RECT 4.975 0.330 6.575 0.490 ;
  END
END XNR2D4

#--------EOF---------

MACRO XOR2D0
  CLASS CORE ;
  FOREIGN XOR2D0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.170300 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 5.600 5.775 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 3.550 4.615 3.680 4.795 ;
        RECT 5.470 4.300 5.600 4.795 ;
        RECT 5.385 4.000 5.685 4.300 ;
        RECT 5.385 2.000 5.685 2.300 ;
        RECT 2.590 1.170 2.720 1.350 ;
        RECT 5.470 1.170 5.600 2.000 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 2.590 0.345 5.600 0.475 ;
      LAYER Metal1 ;
        RECT 5.405 4.070 5.665 4.230 ;
        RECT 5.455 2.230 5.615 4.070 ;
        RECT 5.405 2.070 5.665 2.230 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.124800 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 3.260 4.640 4.600 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 4.425 2.000 4.725 2.300 ;
        RECT 4.510 1.280 4.640 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 4.495 2.230 4.655 3.030 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.542400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 4.615 1.760 4.795 ;
        RECT 0.670 4.215 0.800 4.600 ;
        RECT 2.025 4.215 2.325 4.300 ;
        RECT 0.670 4.085 2.325 4.215 ;
        RECT 2.590 4.215 2.720 4.795 ;
        RECT 2.590 4.085 4.160 4.215 ;
        RECT 0.670 1.280 0.800 4.085 ;
        RECT 2.025 4.000 2.325 4.085 ;
        RECT 4.030 2.695 4.160 4.085 ;
        RECT 5.865 2.695 6.165 2.780 ;
        RECT 4.030 2.565 6.165 2.695 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 1.630 2.085 3.765 2.215 ;
        RECT 1.630 1.170 1.760 2.085 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 4.030 1.555 4.160 2.565 ;
        RECT 5.865 2.480 6.165 2.565 ;
        RECT 3.550 1.425 4.160 1.555 ;
        RECT 3.550 1.170 3.680 1.425 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 3.695 5.790 ;
        RECT 3.535 5.130 3.695 5.630 ;
        RECT 1.615 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 1.615 1.150 1.775 4.970 ;
        RECT 3.055 4.230 3.215 4.970 ;
        RECT 2.045 4.070 3.215 4.230 ;
        RECT 3.055 1.150 3.215 4.070 ;
        RECT 4.015 2.230 4.175 4.970 ;
        RECT 5.935 2.710 6.095 4.970 ;
        RECT 5.885 2.550 6.145 2.710 ;
        RECT 3.485 2.070 4.175 2.230 ;
        RECT 4.015 1.150 4.175 2.070 ;
        RECT 5.935 1.150 6.095 2.550 ;
        RECT 1.615 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
  END
END XOR2D0

#--------EOF---------

MACRO XOR2D1
  CLASS CORE ;
  FOREIGN XOR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 5.600 5.775 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 2.985 3.175 3.285 3.260 ;
        RECT 3.550 3.175 3.680 4.600 ;
        RECT 5.470 4.215 5.600 4.600 ;
        RECT 5.470 4.085 6.080 4.215 ;
        RECT 2.985 3.045 3.680 3.175 ;
        RECT 2.985 2.960 3.285 3.045 ;
        RECT 3.070 1.555 3.200 2.960 ;
        RECT 5.950 2.215 6.080 4.085 ;
        RECT 2.590 1.425 3.200 1.555 ;
        RECT 5.470 2.085 6.080 2.215 ;
        RECT 2.590 1.280 2.720 1.425 ;
        RECT 5.470 1.280 5.600 2.085 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 3.055 3.190 3.215 4.230 ;
        RECT 3.005 3.030 3.265 3.190 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.000 4.725 2.300 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.084800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 0.125 1.410 0.385 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 0.000 -0.150 6.460 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 6.460 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 4.420 1.760 4.600 ;
        RECT 0.670 3.175 0.800 4.000 ;
        RECT 2.025 3.175 2.325 3.260 ;
        RECT 0.670 3.045 2.325 3.175 ;
        RECT 0.670 1.640 0.800 3.045 ;
        RECT 2.025 2.960 2.325 3.045 ;
        RECT 2.590 2.780 2.720 4.600 ;
        RECT 2.505 2.480 2.805 2.780 ;
        RECT 3.465 2.480 3.765 2.780 ;
        RECT 1.630 1.280 1.760 1.460 ;
        RECT 3.550 1.280 3.680 2.480 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 1.545 0.260 1.845 0.560 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 3.695 5.790 ;
        RECT 3.535 5.130 3.695 5.630 ;
        RECT 1.615 4.970 2.305 5.130 ;
        RECT 2.575 4.970 3.265 5.130 ;
        RECT 3.535 4.970 4.225 5.130 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 1.615 1.150 1.775 4.970 ;
        RECT 2.575 3.190 2.735 4.970 ;
        RECT 5.935 4.790 6.095 4.970 ;
        RECT 2.045 3.030 2.735 3.190 ;
        RECT 3.535 4.630 6.095 4.790 ;
        RECT 2.095 2.230 2.255 3.030 ;
        RECT 3.535 2.710 3.695 4.630 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 2.525 2.550 3.745 2.710 ;
        RECT 2.095 2.070 3.215 2.230 ;
        RECT 3.055 1.150 3.215 2.070 ;
        RECT 4.015 1.570 4.175 4.070 ;
        RECT 3.965 1.410 4.225 1.570 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 1.615 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.535 0.990 4.225 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 3.535 0.490 3.695 0.990 ;
        RECT 1.565 0.330 3.695 0.490 ;
  END
END XOR2D1

#--------EOF---------

MACRO XOR2D2
  CLASS CORE ;
  FOREIGN XOR2D2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.645 3.680 5.775 ;
        RECT 0.670 5.200 0.800 5.645 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 0.670 2.695 0.800 4.600 ;
        RECT 3.550 4.420 3.680 4.600 ;
        RECT 2.505 2.695 2.805 2.780 ;
        RECT 0.670 2.565 2.805 2.695 ;
        RECT 0.670 1.280 0.800 2.565 ;
        RECT 2.505 2.480 2.805 2.565 ;
        RECT 2.590 1.280 2.720 2.480 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.095 2.550 2.785 2.710 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249600 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 4.425 2.000 4.725 2.300 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.230 4.655 2.710 ;
        RECT 4.445 2.070 4.705 2.230 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 5.935 1.570 6.095 4.070 ;
        RECT 5.885 1.410 6.145 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 3.175 1.760 4.600 ;
        RECT 2.590 4.215 2.720 4.600 ;
        RECT 2.590 4.085 3.680 4.215 ;
        RECT 2.985 3.175 3.285 3.260 ;
        RECT 1.630 3.045 3.285 3.175 ;
        RECT 2.985 2.960 3.285 3.045 ;
        RECT 2.025 2.000 2.325 2.300 ;
        RECT 2.110 1.555 2.240 2.000 ;
        RECT 1.630 1.425 2.240 1.555 ;
        RECT 1.630 1.280 1.760 1.425 ;
        RECT 3.550 1.280 3.680 4.085 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 3.260 6.560 4.000 ;
        RECT 6.345 2.960 6.645 3.260 ;
        RECT 6.345 2.215 6.645 2.300 ;
        RECT 5.470 2.085 6.645 2.215 ;
        RECT 5.470 1.640 5.600 2.085 ;
        RECT 6.345 2.000 6.645 2.085 ;
        RECT 6.430 1.640 6.560 2.000 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 0.585 0.345 3.680 0.475 ;
        RECT 4.425 0.475 4.725 0.560 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 4.425 0.345 5.600 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
        RECT 4.425 0.260 4.725 0.345 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 2.045 4.970 2.735 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 2.575 3.190 2.735 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 3.055 4.630 6.575 4.790 ;
        RECT 3.965 4.070 4.225 4.230 ;
        RECT 1.615 3.030 2.735 3.190 ;
        RECT 3.005 3.030 3.265 3.190 ;
        RECT 1.615 1.150 1.775 3.030 ;
        RECT 3.055 2.230 3.215 3.030 ;
        RECT 4.015 2.230 4.175 4.070 ;
        RECT 6.415 3.190 6.575 4.630 ;
        RECT 6.365 3.030 6.625 3.190 ;
        RECT 6.415 2.230 6.575 3.030 ;
        RECT 2.045 2.070 4.175 2.230 ;
        RECT 6.365 2.070 6.625 2.230 ;
        RECT 4.015 1.570 4.175 2.070 ;
        RECT 3.965 1.410 4.225 1.570 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 1.615 0.990 2.305 1.150 ;
        RECT 3.005 0.990 4.655 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 4.495 0.490 4.655 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 4.445 0.330 4.705 0.490 ;
  END
END XOR2D2

#--------EOF---------

MACRO XOR2D4
  CLASS CORE ;
  FOREIGN XOR2D4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.713700 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 5.470 2.215 5.600 4.000 ;
        RECT 6.430 2.215 6.560 4.000 ;
        RECT 9.310 2.215 9.440 4.000 ;
        RECT 4.425 2.085 9.440 2.215 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 4.510 1.505 4.640 2.000 ;
        RECT 7.390 1.505 7.520 2.085 ;
        RECT 9.310 1.640 9.440 2.085 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
      LAYER Metal1 ;
        RECT 4.445 2.070 4.705 2.230 ;
        RECT 4.495 1.410 4.655 2.070 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.748800 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 0.670 2.215 0.800 4.000 ;
        RECT 1.630 2.215 1.760 4.000 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 0.670 2.085 2.805 2.215 ;
        RECT 0.670 1.640 0.800 2.085 ;
        RECT 1.630 1.640 1.760 2.085 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.230 2.735 2.710 ;
        RECT 2.525 2.070 2.785 2.230 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.187200 ;
    PORT
      LAYER Metal1 ;
        RECT 10.685 4.070 10.945 4.230 ;
        RECT 12.605 4.070 12.865 4.230 ;
        RECT 10.735 1.570 10.895 4.070 ;
        RECT 12.655 1.570 12.815 4.070 ;
        RECT 10.685 1.410 12.865 1.570 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 9.775 0.150 9.935 0.990 ;
        RECT 11.695 0.150 11.855 0.990 ;
        RECT 13.615 0.150 13.775 0.990 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 9.775 5.130 9.935 5.970 ;
        RECT 11.695 5.130 11.855 5.970 ;
        RECT 13.615 5.130 13.775 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 9.725 4.970 9.985 5.130 ;
        RECT 11.645 4.970 11.905 5.130 ;
        RECT 13.565 4.970 13.825 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 8.265 4.900 8.565 5.200 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 4.510 3.260 4.640 4.000 ;
        RECT 7.390 3.260 7.520 4.000 ;
        RECT 4.425 2.960 4.725 3.260 ;
        RECT 7.305 2.960 7.605 3.260 ;
        RECT 6.825 2.695 7.125 2.780 ;
        RECT 8.350 2.695 8.480 4.900 ;
        RECT 6.825 2.565 8.480 2.695 ;
        RECT 6.825 2.480 7.125 2.565 ;
        RECT 10.270 2.300 10.400 4.000 ;
        RECT 3.465 2.000 3.765 2.300 ;
        RECT 10.185 2.215 10.485 2.300 ;
        RECT 11.230 2.215 11.360 4.000 ;
        RECT 12.190 2.215 12.320 4.000 ;
        RECT 13.150 2.215 13.280 4.000 ;
        RECT 10.185 2.085 13.280 2.215 ;
        RECT 10.185 2.000 10.485 2.085 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 5.470 1.505 5.600 1.685 ;
        RECT 6.430 1.505 6.560 1.685 ;
        RECT 10.270 1.640 10.400 2.000 ;
        RECT 11.230 1.640 11.360 2.085 ;
        RECT 12.190 1.640 12.320 2.085 ;
        RECT 13.150 1.640 13.280 2.085 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 6.430 0.560 6.560 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 6.345 0.475 6.645 0.560 ;
        RECT 5.470 0.345 6.645 0.475 ;
        RECT 6.345 0.260 6.645 0.345 ;
      LAYER Metal1 ;
        RECT 4.015 4.970 8.545 5.130 ;
        RECT 0.125 4.070 0.385 4.230 ;
        RECT 2.045 4.070 2.305 4.230 ;
        RECT 0.175 1.570 0.335 4.070 ;
        RECT 2.095 1.570 2.255 4.070 ;
        RECT 4.015 2.710 4.175 4.970 ;
        RECT 4.495 4.630 6.575 4.790 ;
        RECT 4.495 3.190 4.655 4.630 ;
        RECT 5.885 4.070 6.145 4.230 ;
        RECT 4.445 3.030 4.705 3.190 ;
        RECT 4.015 2.550 5.135 2.710 ;
        RECT 3.485 2.070 3.745 2.230 ;
        RECT 3.535 1.570 3.695 2.070 ;
        RECT 0.125 1.410 3.695 1.570 ;
        RECT 3.535 1.150 3.695 1.410 ;
        RECT 4.975 1.150 5.135 2.550 ;
        RECT 5.935 1.150 6.095 4.070 ;
        RECT 6.415 3.190 6.575 4.630 ;
        RECT 8.765 4.070 9.025 4.230 ;
        RECT 8.815 3.190 8.975 4.070 ;
        RECT 6.415 3.030 8.975 3.190 ;
        RECT 3.535 0.990 6.145 1.150 ;
        RECT 6.415 0.490 6.575 3.030 ;
        RECT 6.845 2.550 7.105 2.710 ;
        RECT 6.895 2.230 7.055 2.550 ;
        RECT 6.895 2.070 10.465 2.230 ;
        RECT 6.895 1.150 7.055 2.070 ;
        RECT 6.845 0.990 9.025 1.150 ;
        RECT 6.895 0.490 7.055 0.990 ;
        RECT 6.365 0.330 7.055 0.490 ;
  END
END XOR2D4

#--------EOF---------


END LIBRARY
