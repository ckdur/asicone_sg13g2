VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SARADC_FILLTIE2
  CLASS BLOCK ;
  FOREIGN SARADC_FILLTIE2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.380 BY 6.120 ;
  SYMMETRY X Y R90 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.590 0.920 0.850 1.080 ;
        RECT 1.070 0.920 1.330 1.080 ;
        RECT 1.550 0.920 1.810 1.080 ;
        RECT 0.640 0.150 0.800 0.920 ;
        RECT 1.120 0.150 1.280 0.920 ;
        RECT 1.600 0.150 1.760 0.920 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.380 6.270 ;
        RECT 0.640 5.200 0.800 5.970 ;
        RECT 1.120 5.200 1.280 5.970 ;
        RECT 1.600 5.200 1.760 5.970 ;
        RECT 0.590 5.040 0.850 5.200 ;
        RECT 1.070 5.040 1.330 5.200 ;
        RECT 1.550 5.040 1.810 5.200 ;
    END
  END vdd
END SARADC_FILLTIE2
END LIBRARY

