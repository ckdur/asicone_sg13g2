VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SARADC_CELL_INVX0_ASSW
  CLASS BLOCK ;
  FOREIGN SARADC_CELL_INVX0_ASSW ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  PIN zn
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN i
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.300 0.800 4.600 ;
        RECT 0.585 2.000 0.885 2.300 ;
        RECT 0.670 1.280 0.800 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.230 0.815 2.710 ;
        RECT 0.605 2.070 0.865 2.230 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 0.175 5.130 0.335 5.970 ;
        RECT 0.125 4.970 0.385 5.130 ;
    END
  END vdd
END SARADC_CELL_INVX0_ASSW
END LIBRARY

