VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SARADC_CELL_INVX16_ASCAP
  CLASS BLOCK ;
  FOREIGN SARADC_CELL_INVX16_ASCAP ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.980 BY 6.120 ;
  SYMMETRY X Y R90 ;
  PIN i
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 0.670 2.300 0.800 4.000 ;
        RECT 1.630 2.300 1.760 4.000 ;
        RECT 2.590 2.300 2.720 4.000 ;
        RECT 3.550 2.300 3.680 4.000 ;
        RECT 4.510 2.300 4.640 4.000 ;
        RECT 5.470 2.300 5.600 4.000 ;
        RECT 6.430 2.300 6.560 4.000 ;
        RECT 7.390 2.300 7.520 4.000 ;
        RECT 8.350 2.300 8.480 4.000 ;
        RECT 9.310 2.300 9.440 4.000 ;
        RECT 10.270 2.300 10.400 4.000 ;
        RECT 11.230 2.300 11.360 4.000 ;
        RECT 12.190 2.300 12.320 4.000 ;
        RECT 13.150 2.300 13.280 4.000 ;
        RECT 14.110 2.300 14.240 4.000 ;
        RECT 15.070 2.300 15.200 4.000 ;
        RECT 0.585 2.215 0.885 2.300 ;
        RECT 1.545 2.215 1.845 2.300 ;
        RECT 2.505 2.215 2.805 2.300 ;
        RECT 3.465 2.215 3.765 2.300 ;
        RECT 4.425 2.215 4.725 2.300 ;
        RECT 5.385 2.215 5.685 2.300 ;
        RECT 6.345 2.215 6.645 2.300 ;
        RECT 7.305 2.215 7.605 2.300 ;
        RECT 8.265 2.215 8.565 2.300 ;
        RECT 9.225 2.215 9.525 2.300 ;
        RECT 10.185 2.215 10.485 2.300 ;
        RECT 11.145 2.215 11.445 2.300 ;
        RECT 12.105 2.215 12.405 2.300 ;
        RECT 13.065 2.215 13.365 2.300 ;
        RECT 14.025 2.215 14.325 2.300 ;
        RECT 14.985 2.215 15.285 2.300 ;
        RECT 0.585 2.085 15.285 2.215 ;
        RECT 0.585 2.000 0.885 2.085 ;
        RECT 1.545 2.000 1.845 2.085 ;
        RECT 2.505 2.000 2.805 2.085 ;
        RECT 3.465 2.000 3.765 2.085 ;
        RECT 4.425 2.000 4.725 2.085 ;
        RECT 5.385 2.000 5.685 2.085 ;
        RECT 6.345 2.000 6.645 2.085 ;
        RECT 7.305 2.000 7.605 2.085 ;
        RECT 8.265 2.000 8.565 2.085 ;
        RECT 9.225 2.000 9.525 2.085 ;
        RECT 10.185 2.000 10.485 2.085 ;
        RECT 11.145 2.000 11.445 2.085 ;
        RECT 12.105 2.000 12.405 2.085 ;
        RECT 13.065 2.000 13.365 2.085 ;
        RECT 14.025 2.000 14.325 2.085 ;
        RECT 14.985 2.000 15.285 2.085 ;
        RECT 0.670 1.640 0.800 2.000 ;
        RECT 1.630 1.640 1.760 2.000 ;
        RECT 2.590 1.640 2.720 2.000 ;
        RECT 3.550 1.640 3.680 2.000 ;
        RECT 4.510 1.640 4.640 2.000 ;
        RECT 5.470 1.640 5.600 2.000 ;
        RECT 6.430 1.640 6.560 2.000 ;
        RECT 7.390 1.640 7.520 2.000 ;
        RECT 8.350 1.640 8.480 2.000 ;
        RECT 9.310 1.640 9.440 2.000 ;
        RECT 10.270 1.640 10.400 2.000 ;
        RECT 11.230 1.640 11.360 2.000 ;
        RECT 12.190 1.640 12.320 2.000 ;
        RECT 13.150 1.640 13.280 2.000 ;
        RECT 14.110 1.640 14.240 2.000 ;
        RECT 15.070 1.640 15.200 2.000 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 15.070 0.740 15.200 0.920 ;
      LAYER Metal1 ;
        RECT 0.605 2.070 15.265 2.230 ;
    END
  END i
  PIN zn
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.070 15.745 4.230 ;
        RECT 15.535 1.570 15.695 4.070 ;
        RECT 0.125 1.410 15.745 1.570 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 12.655 0.150 12.815 0.990 ;
        RECT 14.575 0.150 14.735 0.990 ;
        RECT 0.000 -0.150 15.980 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 15.980 6.270 ;
        RECT 1.135 5.130 1.295 5.970 ;
        RECT 3.055 5.130 3.215 5.970 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 6.895 5.130 7.055 5.970 ;
        RECT 8.815 5.130 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 12.655 5.130 12.815 5.970 ;
        RECT 14.575 5.130 14.735 5.970 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 14.525 4.970 14.785 5.130 ;
    END
  END vdd
END SARADC_CELL_INVX16_ASCAP
END LIBRARY

