VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.34 BY 6.12 ;
END obssite

#--------EOF---------

MACRO AN2D1
  CLASS CORE ;
  FOREIGN AN2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.025 3.635 2.325 3.720 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 2.025 3.505 3.680 3.635 ;
        RECT 2.025 3.420 2.325 3.505 ;
        RECT 3.550 1.620 3.680 3.505 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.630 1.775 4.790 ;
        RECT 1.615 3.650 1.775 4.630 ;
        RECT 1.615 3.490 2.305 3.650 ;
        RECT 2.095 1.150 2.255 3.490 ;
        RECT 2.045 0.990 2.305 1.150 ;
  END
END AN2D1

#--------EOF---------

MACRO AN2D1_1
  CLASS CORE ;
  FOREIGN AN2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 1.390 0.815 2.050 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.050 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.760 2.720 4.100 ;
        RECT 2.505 2.460 2.805 2.760 ;
        RECT 2.590 1.620 2.720 2.460 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 2.690 1.295 4.630 ;
        RECT 0.175 2.530 2.785 2.690 ;
        RECT 0.175 1.150 0.335 2.530 ;
        RECT 0.125 0.990 0.385 1.150 ;
  END
END AN2D1_1

#--------EOF---------

MACRO AN2D1_2
  CLASS CORE ;
  FOREIGN AN2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.025 3.635 2.325 3.720 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 2.025 3.505 3.680 3.635 ;
        RECT 2.025 3.420 2.325 3.505 ;
        RECT 3.550 1.620 3.680 3.505 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 2.095 3.650 2.255 4.630 ;
        RECT 0.655 3.490 2.305 3.650 ;
        RECT 2.095 1.150 2.255 3.490 ;
        RECT 2.045 0.990 2.305 1.150 ;
  END
END AN2D1_2

#--------EOF---------

MACRO AN2D1_3
  CLASS CORE ;
  FOREIGN AN2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.025 3.635 2.325 3.720 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 2.025 3.505 3.680 3.635 ;
        RECT 2.025 3.420 2.325 3.505 ;
        RECT 3.550 1.620 3.680 3.505 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 2.305 4.790 ;
        RECT 2.095 3.650 2.255 4.630 ;
        RECT 2.045 3.490 2.305 3.650 ;
        RECT 2.095 1.150 2.255 3.490 ;
        RECT 0.125 0.990 2.255 1.150 ;
  END
END AN2D1_3

#--------EOF---------

MACRO AO21D1
  CLASS CORE ;
  FOREIGN AO21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.545 2.460 1.845 2.760 ;
        RECT 1.630 1.620 1.760 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 1.615 2.690 1.775 3.490 ;
        RECT 1.565 2.530 1.825 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 3.720 2.720 4.100 ;
        RECT 2.505 3.420 2.805 3.720 ;
        RECT 2.505 2.460 2.805 2.760 ;
        RECT 2.590 1.620 2.720 2.460 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 3.490 2.785 3.650 ;
        RECT 2.575 2.690 2.735 3.490 ;
        RECT 2.525 2.530 2.785 2.690 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 1.150 4.175 4.630 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.065 3.155 1.365 3.240 ;
        RECT 2.985 3.155 3.285 3.240 ;
        RECT 4.510 3.155 4.640 4.100 ;
        RECT 1.065 3.025 4.640 3.155 ;
        RECT 1.065 2.940 1.365 3.025 ;
        RECT 2.985 2.940 3.285 3.025 ;
        RECT 4.510 1.620 4.640 1.800 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 2.985 0.345 4.640 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.330 0.335 4.630 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 3.055 3.170 3.215 4.970 ;
        RECT 1.085 3.010 1.345 3.170 ;
        RECT 3.005 3.010 3.265 3.170 ;
        RECT 1.135 1.150 1.295 3.010 ;
        RECT 3.055 1.150 3.215 3.010 ;
        RECT 0.125 0.990 1.295 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END AO21D1

#--------EOF---------

MACRO AO21D1_1
  CLASS CORE ;
  FOREIGN AO21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 1.150 5.135 4.630 ;
        RECT 4.925 0.990 5.185 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.505 4.560 2.805 4.860 ;
        RECT 2.590 3.720 2.720 4.560 ;
        RECT 4.510 3.720 4.640 4.100 ;
        RECT 2.505 3.420 2.805 3.720 ;
        RECT 4.425 3.420 4.725 3.720 ;
        RECT 2.590 1.220 2.720 3.420 ;
        RECT 4.510 1.620 4.640 3.420 ;
        RECT 2.505 0.920 2.805 1.220 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.045 4.630 2.785 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 2.525 3.490 4.705 3.650 ;
        RECT 2.045 0.990 3.265 1.150 ;
  END
END AO21D1_1

#--------EOF---------

MACRO AO21D1_2
  CLASS CORE ;
  FOREIGN AO21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.630 4.655 4.790 ;
        RECT 4.495 1.150 4.655 4.630 ;
        RECT 3.965 0.990 4.655 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 3.945 3.635 4.245 3.720 ;
        RECT 4.510 3.635 4.640 4.100 ;
        RECT 3.945 3.505 4.640 3.635 ;
        RECT 3.945 3.420 4.245 3.505 ;
        RECT 4.510 1.620 4.640 1.800 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.260 4.725 0.560 ;
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 1.135 1.150 1.295 4.170 ;
        RECT 4.015 3.650 4.175 4.170 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 1.135 0.330 4.705 0.490 ;
  END
END AO21D1_2

#--------EOF---------

MACRO AO21D1_3
  CLASS CORE ;
  FOREIGN AO21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 1.150 4.175 4.630 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 1.620 4.640 4.100 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 2.985 0.345 4.640 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 2.095 4.170 3.215 4.330 ;
        RECT 3.055 1.150 3.215 4.170 ;
        RECT 0.125 0.990 3.265 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 3.005 0.330 3.265 0.490 ;
  END
END AO21D1_3

#--------EOF---------

MACRO AOI21D1
  CLASS CORE ;
  FOREIGN AOI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.494000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 1.150 2.255 4.170 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 3.055 4.790 3.215 5.970 ;
        RECT 3.005 4.630 3.265 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
  END
END AOI21D1

#--------EOF---------

MACRO AOI21D1_1
  CLASS CORE ;
  FOREIGN AOI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.494000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 1.150 1.295 4.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
  END
END AOI21D1_1

#--------EOF---------

MACRO AOI21D1_2
  CLASS CORE ;
  FOREIGN AOI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.034000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.655 4.330 0.815 4.630 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 0.655 4.170 2.255 4.330 ;
        RECT 0.655 1.150 0.815 4.170 ;
        RECT 0.655 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.105 2.195 0.405 2.280 ;
        RECT 0.670 2.195 0.800 4.100 ;
        RECT 0.105 2.065 0.800 2.195 ;
        RECT 0.105 1.980 0.405 2.065 ;
        RECT 0.670 1.620 0.800 2.065 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 2.210 0.335 2.690 ;
        RECT 0.125 2.050 0.385 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
  END
END AOI21D1_2

#--------EOF---------

MACRO AOI21D1_3
  CLASS CORE ;
  FOREIGN AOI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.034000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.330 0.335 4.630 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 2.095 1.150 2.255 4.170 ;
        RECT 0.125 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.790 1.295 4.970 ;
        RECT 3.055 4.790 3.215 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
  END
END AOI21D1_3

#--------EOF---------

MACRO ANTENNA
  CLASS CORE ANTENNACELL ;
  FOREIGN ANTENNA ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.380 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.380 6.270 ;
    END
  END vdd
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.440450 ;
    ANTENNADIFFAREA 2.880900 ;
    PORT
      LAYER Metal1 ;
        RECT 0.590 5.040 1.810 5.200 ;
        RECT 0.640 1.080 0.800 5.040 ;
        RECT 0.590 0.920 1.810 1.080 ;
    END
  END i
END ANTENNA

#--------EOF---------

MACRO BUFFD1
  CLASS CORE ;
  FOREIGN BUFFD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.650 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.270 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.670 2.280 0.800 3.420 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 4.970 2.305 5.130 ;
        RECT 1.615 3.650 1.775 4.970 ;
        RECT 0.605 3.490 1.775 3.650 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 1.150 0.815 2.050 ;
        RECT 0.655 0.990 2.305 1.150 ;
  END
END BUFFD1

#--------EOF---------

MACRO BUFFD1_1
  CLASS CORE ;
  FOREIGN BUFFD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.650 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.270 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.630 2.280 1.760 3.420 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 0.655 3.650 0.815 4.970 ;
        RECT 0.655 3.490 1.825 3.650 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.150 1.775 2.050 ;
        RECT 0.125 0.990 1.775 1.150 ;
  END
END BUFFD1_1

#--------EOF---------

MACRO BUFFD1_2
  CLASS CORE ;
  FOREIGN BUFFD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.650 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.270 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.630 2.280 1.760 3.420 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 0.655 3.650 0.815 4.970 ;
        RECT 0.655 3.490 1.825 3.650 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.150 1.775 2.050 ;
        RECT 0.125 0.990 1.775 1.150 ;
  END
END BUFFD1_2

#--------EOF---------

MACRO BUFFD1_3
  CLASS CORE ;
  FOREIGN BUFFD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.650 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.270 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.630 2.280 1.760 3.420 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 0.655 3.650 0.815 4.970 ;
        RECT 0.655 3.490 1.825 3.650 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.150 1.775 2.050 ;
        RECT 0.125 0.990 1.775 1.150 ;
  END
END BUFFD1_3

#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ;
  FOREIGN DFCNQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.000 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.117000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.155 0.800 4.650 ;
        RECT 0.190 3.025 0.800 3.155 ;
        RECT 0.190 2.280 0.320 3.025 ;
        RECT 0.105 1.980 0.405 2.280 ;
        RECT 0.190 1.535 0.320 1.980 ;
        RECT 0.190 1.405 0.800 1.535 ;
        RECT 0.670 1.270 0.800 1.405 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 2.210 0.335 2.690 ;
        RECT 0.125 2.050 0.385 2.210 ;
    END
  END cp
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150800 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.390 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.270 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 1.390 4.655 2.050 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.287300 ;
    PORT
      LAYER GatPoly ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 8.350 4.775 8.480 4.925 ;
        RECT 7.390 4.645 8.480 4.775 ;
        RECT 7.390 1.620 7.520 4.645 ;
        RECT 13.150 3.720 13.280 4.210 ;
        RECT 13.065 3.420 13.365 3.720 ;
        RECT 13.065 1.980 13.365 2.280 ;
        RECT 13.150 1.620 13.280 1.980 ;
        RECT 7.305 1.320 7.605 1.620 ;
        RECT 7.390 1.165 7.520 1.320 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 13.150 0.740 13.280 0.920 ;
      LAYER Metal1 ;
        RECT 13.085 3.490 13.345 3.650 ;
        RECT 13.135 2.210 13.295 3.490 ;
        RECT 11.215 2.050 13.345 2.210 ;
        RECT 11.215 1.550 11.375 2.050 ;
        RECT 7.325 1.390 11.375 1.550 ;
    END
  END cdn
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.485 4.630 16.655 4.790 ;
        RECT 16.495 1.150 16.655 4.630 ;
        RECT 16.445 0.990 16.705 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 17.000 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 5.385 5.560 5.685 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.560 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 14.110 5.200 14.240 5.380 ;
        RECT 15.070 5.200 15.200 5.380 ;
        RECT 5.470 4.690 5.600 4.870 ;
        RECT 1.630 2.760 1.760 4.650 ;
        RECT 3.550 3.720 3.680 4.390 ;
        RECT 6.430 3.720 6.560 4.895 ;
        RECT 3.465 3.420 3.765 3.720 ;
        RECT 6.345 3.420 6.645 3.720 ;
        RECT 0.585 2.675 0.885 2.760 ;
        RECT 1.545 2.675 1.845 2.760 ;
        RECT 0.585 2.545 1.845 2.675 ;
        RECT 0.585 2.460 0.885 2.545 ;
        RECT 1.545 2.460 1.845 2.545 ;
        RECT 1.630 1.270 1.760 2.460 ;
        RECT 3.550 2.280 3.680 3.420 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 6.430 1.620 6.560 3.420 ;
        RECT 8.265 2.940 8.565 3.240 ;
        RECT 8.350 2.280 8.480 2.940 ;
        RECT 9.310 2.280 9.440 4.485 ;
        RECT 10.270 2.760 10.400 4.170 ;
        RECT 10.185 2.460 10.485 2.760 ;
        RECT 8.265 1.980 8.565 2.280 ;
        RECT 9.225 1.980 9.525 2.280 ;
        RECT 2.505 1.535 2.805 1.620 ;
        RECT 2.505 1.405 3.680 1.535 ;
        RECT 2.505 1.320 2.805 1.405 ;
        RECT 3.550 1.270 3.680 1.405 ;
        RECT 5.470 1.165 5.600 1.345 ;
        RECT 6.345 1.320 6.645 1.620 ;
        RECT 8.350 1.350 8.480 1.980 ;
        RECT 9.310 1.410 9.440 1.590 ;
        RECT 6.430 1.165 6.560 1.320 ;
        RECT 10.270 1.165 10.400 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 5.470 0.560 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.560 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 5.385 0.260 5.685 0.560 ;
        RECT 9.225 0.475 9.525 0.560 ;
        RECT 11.230 0.475 11.360 4.925 ;
        RECT 12.190 3.155 12.320 4.925 ;
        RECT 14.110 3.720 14.240 4.210 ;
        RECT 14.025 3.420 14.325 3.720 ;
        RECT 13.545 3.155 13.845 3.240 ;
        RECT 15.070 3.155 15.200 4.100 ;
        RECT 12.190 3.025 16.160 3.155 ;
        RECT 12.190 1.620 12.320 3.025 ;
        RECT 13.545 2.940 13.845 3.025 ;
        RECT 14.025 2.460 14.325 2.760 ;
        RECT 14.110 1.620 14.240 2.460 ;
        RECT 16.030 1.620 16.160 3.025 ;
        RECT 12.105 1.320 12.405 1.620 ;
        RECT 12.190 1.165 12.320 1.320 ;
        RECT 12.190 0.740 12.320 0.920 ;
        RECT 14.110 0.560 14.240 0.920 ;
        RECT 16.030 0.740 16.160 0.920 ;
        RECT 9.225 0.345 11.360 0.475 ;
        RECT 9.225 0.260 9.525 0.345 ;
        RECT 14.025 0.260 14.325 0.560 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 5.665 5.790 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 2.045 4.970 3.695 5.130 ;
        RECT 5.885 4.970 8.065 5.130 ;
        RECT 10.685 4.970 14.255 5.130 ;
        RECT 0.655 2.690 0.815 4.970 ;
        RECT 3.535 3.650 3.695 4.970 ;
        RECT 4.925 4.630 5.615 4.790 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 5.455 3.170 5.615 4.630 ;
        RECT 9.295 4.630 9.985 4.790 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 9.295 3.650 9.455 4.630 ;
        RECT 6.365 3.490 9.455 3.650 ;
        RECT 13.615 3.170 13.775 4.630 ;
        RECT 14.095 3.650 14.255 4.970 ;
        RECT 14.045 3.490 14.305 3.650 ;
        RECT 5.455 3.010 8.545 3.170 ;
        RECT 13.565 3.010 13.825 3.170 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 2.575 2.530 10.465 2.690 ;
        RECT 1.615 1.550 1.775 2.530 ;
        RECT 2.575 1.550 2.735 2.530 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 4.975 2.050 9.505 2.210 ;
        RECT 0.175 1.390 2.785 1.550 ;
        RECT 0.175 1.150 0.335 1.390 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 3.535 0.490 3.695 2.050 ;
        RECT 4.975 1.150 5.135 2.050 ;
        RECT 13.615 1.550 13.775 3.010 ;
        RECT 14.095 2.690 14.255 3.490 ;
        RECT 14.045 2.530 14.305 2.690 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 12.125 1.390 14.735 1.550 ;
        RECT 6.415 1.150 6.575 1.390 ;
        RECT 14.575 1.150 14.735 1.390 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.415 0.990 9.025 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 10.685 0.990 11.905 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 9.775 0.490 9.935 0.990 ;
        RECT 2.095 0.330 9.505 0.490 ;
        RECT 9.775 0.330 14.305 0.490 ;
  END
END DFCNQD1

#--------EOF---------

MACRO DFQD1
  CLASS CORE ;
  FOREIGN DFQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.960 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.142350 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 4.400 2.720 4.510 ;
        RECT 2.505 4.100 2.805 4.400 ;
        RECT 2.590 1.325 2.720 1.505 ;
        RECT 2.590 0.560 2.720 0.920 ;
        RECT 2.505 0.260 2.805 0.560 ;
      LAYER Metal1 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 2.575 0.490 2.735 4.170 ;
        RECT 2.525 0.330 2.785 0.490 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.585 2.460 0.885 2.760 ;
        RECT 0.670 1.620 0.800 2.460 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 2.690 0.815 3.490 ;
        RECT 0.605 2.530 0.865 2.690 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 13.615 1.150 13.775 4.630 ;
        RECT 13.565 0.990 13.825 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 8.815 0.150 8.975 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 14.960 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.960 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 8.815 4.790 8.975 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.105 5.775 0.405 5.860 ;
        RECT 3.465 5.775 3.765 5.860 ;
        RECT 0.105 5.645 3.765 5.775 ;
        RECT 0.105 5.560 0.405 5.645 ;
        RECT 3.465 5.560 3.765 5.645 ;
        RECT 5.385 5.775 5.685 5.860 ;
        RECT 5.385 5.645 7.520 5.775 ;
        RECT 5.385 5.560 5.685 5.645 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.560 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 5.470 5.200 5.600 5.560 ;
        RECT 7.390 5.200 7.520 5.645 ;
        RECT 11.230 5.645 14.240 5.775 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 11.230 5.200 11.360 5.645 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 14.110 5.200 14.240 5.645 ;
        RECT 3.550 4.745 3.680 4.925 ;
        RECT 1.630 3.635 1.760 4.390 ;
        RECT 3.465 4.100 3.765 4.400 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 1.630 3.505 3.680 3.635 ;
        RECT 0.105 3.155 0.405 3.240 ;
        RECT 0.105 3.025 1.760 3.155 ;
        RECT 0.105 2.940 0.405 3.025 ;
        RECT 1.630 1.325 1.760 3.025 ;
        RECT 3.550 1.165 3.680 3.505 ;
        RECT 4.510 1.165 4.640 4.925 ;
        RECT 8.350 4.400 8.480 4.510 ;
        RECT 11.230 4.400 11.360 4.925 ;
        RECT 5.470 1.620 5.600 4.100 ;
        RECT 7.390 4.045 7.520 4.225 ;
        RECT 8.265 4.100 8.565 4.400 ;
        RECT 11.145 4.100 11.445 4.400 ;
        RECT 9.310 3.720 9.440 4.100 ;
        RECT 9.225 3.420 9.525 3.720 ;
        RECT 6.825 3.155 7.125 3.240 ;
        RECT 9.310 3.155 9.440 3.420 ;
        RECT 11.230 3.240 11.360 4.100 ;
        RECT 6.825 3.025 9.440 3.155 ;
        RECT 6.825 2.940 7.125 3.025 ;
        RECT 11.145 2.940 11.445 3.240 ;
        RECT 12.190 2.675 12.320 4.925 ;
        RECT 12.585 3.420 12.885 3.720 ;
        RECT 7.390 2.545 12.320 2.675 ;
        RECT 6.345 1.535 6.645 1.620 ;
        RECT 7.390 1.535 7.520 2.545 ;
        RECT 8.265 1.980 8.565 2.280 ;
        RECT 12.670 2.195 12.800 3.420 ;
        RECT 9.310 2.065 12.800 2.195 ;
        RECT 6.345 1.405 7.520 1.535 ;
        RECT 6.345 1.320 6.645 1.405 ;
        RECT 7.390 1.295 7.520 1.405 ;
        RECT 8.350 1.375 8.480 1.980 ;
        RECT 9.310 1.620 9.440 2.065 ;
        RECT 14.110 1.620 14.240 4.100 ;
        RECT 11.145 1.320 11.445 1.620 ;
        RECT 11.230 1.165 11.360 1.320 ;
        RECT 12.190 1.165 12.320 1.345 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.260 4.725 0.560 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 12.190 0.475 12.320 0.920 ;
        RECT 14.110 0.740 14.240 0.920 ;
        RECT 5.470 0.345 12.320 0.475 ;
      LAYER Metal1 ;
        RECT 0.125 5.630 0.385 5.790 ;
        RECT 3.485 5.630 5.665 5.790 ;
        RECT 0.175 4.790 0.335 5.630 ;
        RECT 3.005 4.970 8.495 5.130 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 0.175 3.170 0.335 4.630 ;
        RECT 0.125 3.010 0.385 3.170 ;
        RECT 0.175 1.150 0.335 3.010 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 5.935 4.330 6.095 4.630 ;
        RECT 3.485 4.170 6.095 4.330 ;
        RECT 5.935 1.550 6.095 4.170 ;
        RECT 6.895 3.170 7.055 4.630 ;
        RECT 6.845 3.010 7.105 3.170 ;
        RECT 5.935 1.390 6.625 1.550 ;
        RECT 5.935 1.150 6.095 1.390 ;
        RECT 6.895 1.150 7.055 3.010 ;
        RECT 7.855 1.150 8.015 4.630 ;
        RECT 8.335 4.330 8.495 4.970 ;
        RECT 9.725 4.630 11.375 4.790 ;
        RECT 11.215 4.330 11.375 4.630 ;
        RECT 8.285 4.170 8.545 4.330 ;
        RECT 11.165 4.170 11.425 4.330 ;
        RECT 8.335 2.210 8.495 4.170 ;
        RECT 12.655 3.650 12.815 4.970 ;
        RECT 9.245 3.490 12.865 3.650 ;
        RECT 11.165 3.010 11.425 3.170 ;
        RECT 8.285 2.050 8.545 2.210 ;
        RECT 11.215 1.550 11.375 3.010 ;
        RECT 9.775 1.390 11.425 1.550 ;
        RECT 9.775 1.150 9.935 1.390 ;
        RECT 12.655 1.150 12.815 3.490 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 7.855 0.490 8.015 0.990 ;
        RECT 4.445 0.330 8.015 0.490 ;
  END
END DFQD1

#--------EOF---------

MACRO DFQD1_1
  CLASS CORE ;
  FOREIGN DFQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.142350 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 4.400 2.720 4.510 ;
        RECT 2.505 4.100 2.805 4.400 ;
        RECT 2.505 2.940 2.805 3.240 ;
        RECT 2.590 1.325 2.720 2.940 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 2.575 3.170 2.735 4.170 ;
        RECT 2.525 3.010 2.785 3.170 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 1.150 12.815 4.630 ;
        RECT 12.605 0.990 12.865 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 4.975 0.150 5.135 0.990 ;
        RECT 6.895 0.150 7.055 0.990 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
        RECT 4.975 5.130 5.135 5.970 ;
        RECT 4.925 4.970 5.185 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.465 5.560 3.765 5.860 ;
        RECT 4.510 5.645 6.560 5.775 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.560 ;
        RECT 4.510 5.200 4.640 5.645 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 3.550 4.745 3.680 4.925 ;
        RECT 4.510 4.745 4.640 4.925 ;
        RECT 6.430 4.860 6.560 5.645 ;
        RECT 9.225 5.560 9.525 5.860 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.560 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 6.345 4.560 6.645 4.860 ;
        RECT 7.390 4.400 7.520 4.510 ;
        RECT 1.630 3.635 1.760 4.390 ;
        RECT 3.465 4.100 3.765 4.400 ;
        RECT 7.305 4.100 7.605 4.400 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 1.630 3.505 3.680 3.635 ;
        RECT 1.545 2.940 1.845 3.240 ;
        RECT 1.630 1.325 1.760 2.940 ;
        RECT 3.550 1.165 3.680 3.505 ;
        RECT 5.470 3.635 5.600 4.100 ;
        RECT 8.350 3.635 8.480 4.225 ;
        RECT 5.470 3.505 8.480 3.635 ;
        RECT 5.470 1.620 5.600 3.505 ;
        RECT 8.350 2.760 8.480 3.505 ;
        RECT 9.310 3.155 9.440 4.925 ;
        RECT 8.830 3.025 9.440 3.155 ;
        RECT 8.265 2.460 8.565 2.760 ;
        RECT 7.305 1.980 7.605 2.280 ;
        RECT 8.830 2.195 8.960 3.025 ;
        RECT 9.225 2.460 9.525 2.760 ;
        RECT 8.350 2.065 8.960 2.195 ;
        RECT 4.425 1.320 4.725 1.620 ;
        RECT 7.390 1.375 7.520 1.980 ;
        RECT 4.510 1.165 4.640 1.320 ;
        RECT 8.350 1.295 8.480 2.065 ;
        RECT 9.310 1.165 9.440 2.460 ;
        RECT 10.270 1.165 10.400 4.925 ;
        RECT 12.105 4.560 12.405 4.860 ;
        RECT 11.230 2.280 11.360 4.100 ;
        RECT 12.190 3.635 12.320 4.560 ;
        RECT 13.150 3.635 13.280 4.100 ;
        RECT 12.190 3.505 13.280 3.635 ;
        RECT 11.145 1.980 11.445 2.280 ;
        RECT 11.230 1.620 11.360 1.980 ;
        RECT 13.150 1.620 13.280 3.505 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 1.630 0.345 5.600 0.475 ;
        RECT 5.865 0.475 6.165 0.560 ;
        RECT 8.350 0.475 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 5.865 0.345 8.480 0.475 ;
        RECT 10.270 0.475 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 11.625 0.475 11.925 0.560 ;
        RECT 13.150 0.475 13.280 0.920 ;
        RECT 10.270 0.345 13.280 0.475 ;
        RECT 5.865 0.260 6.165 0.345 ;
        RECT 11.625 0.260 11.925 0.345 ;
      LAYER Metal1 ;
        RECT 0.655 5.630 3.745 5.790 ;
        RECT 5.935 5.630 9.505 5.790 ;
        RECT 0.655 4.790 0.815 5.630 ;
        RECT 5.935 4.790 6.095 5.630 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 6.365 4.630 8.065 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 11.645 4.630 12.385 4.790 ;
        RECT 0.655 3.170 0.815 4.630 ;
        RECT 3.055 3.170 3.215 4.630 ;
        RECT 5.935 4.330 6.095 4.630 ;
        RECT 3.485 4.170 6.095 4.330 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 7.375 3.170 7.535 4.170 ;
        RECT 0.175 3.010 1.825 3.170 ;
        RECT 3.055 3.010 7.535 3.170 ;
        RECT 0.175 1.150 0.335 3.010 ;
        RECT 3.055 2.210 3.215 3.010 ;
        RECT 3.055 2.050 7.585 2.210 ;
        RECT 3.055 1.150 3.215 2.050 ;
        RECT 7.855 1.550 8.015 4.630 ;
        RECT 8.815 4.330 8.975 4.630 ;
        RECT 8.815 4.170 9.935 4.330 ;
        RECT 8.285 2.530 9.505 2.690 ;
        RECT 9.775 2.210 9.935 4.170 ;
        RECT 4.445 1.390 8.015 1.550 ;
        RECT 7.855 1.150 8.015 1.390 ;
        RECT 8.815 2.050 11.425 2.210 ;
        RECT 8.815 1.150 8.975 2.050 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 5.935 0.490 6.095 0.990 ;
        RECT 11.695 0.490 11.855 0.990 ;
        RECT 5.885 0.330 6.145 0.490 ;
        RECT 11.645 0.330 11.905 0.490 ;
  END
END DFQD1_1

#--------EOF---------

MACRO DFQD1_2
  CLASS CORE ;
  FOREIGN DFQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.142350 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.510 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.325 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 1.150 12.815 4.630 ;
        RECT 12.605 0.990 12.865 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 8.265 5.775 8.565 5.860 ;
        RECT 8.265 5.645 9.440 5.775 ;
        RECT 8.265 5.560 8.565 5.645 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.645 ;
        RECT 11.145 5.560 11.445 5.860 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.560 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 2.505 4.560 2.805 4.860 ;
        RECT 2.590 4.315 2.720 4.560 ;
        RECT 3.550 4.315 3.680 4.390 ;
        RECT 2.590 4.185 3.680 4.315 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.630 2.280 1.760 3.420 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 2.590 0.560 2.720 4.185 ;
        RECT 4.905 4.100 5.205 4.400 ;
        RECT 4.990 2.760 5.120 4.100 ;
        RECT 5.470 3.720 5.600 4.925 ;
        RECT 6.430 4.400 6.560 4.925 ;
        RECT 9.310 4.745 9.440 4.925 ;
        RECT 6.345 4.100 6.645 4.400 ;
        RECT 5.385 3.420 5.685 3.720 ;
        RECT 4.905 2.460 5.205 2.760 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.325 3.680 1.980 ;
        RECT 6.430 1.620 6.560 4.100 ;
        RECT 7.390 2.760 7.520 4.510 ;
        RECT 8.350 3.720 8.480 4.225 ;
        RECT 8.265 3.635 8.565 3.720 ;
        RECT 8.265 3.505 9.440 3.635 ;
        RECT 8.265 3.420 8.565 3.505 ;
        RECT 7.305 2.460 7.605 2.760 ;
        RECT 5.470 1.165 5.600 1.345 ;
        RECT 6.345 1.320 6.645 1.620 ;
        RECT 7.390 1.375 7.520 2.460 ;
        RECT 6.430 1.165 6.560 1.320 ;
        RECT 8.350 1.295 8.480 1.475 ;
        RECT 9.310 1.165 9.440 3.505 ;
        RECT 10.270 1.620 10.400 4.925 ;
        RECT 11.230 3.920 11.360 4.100 ;
        RECT 11.230 1.620 11.360 1.800 ;
        RECT 13.150 1.620 13.280 4.100 ;
        RECT 10.185 1.320 10.485 1.620 ;
        RECT 10.270 1.165 10.400 1.320 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 5.470 0.560 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.560 8.480 0.920 ;
        RECT 9.310 0.740 9.440 0.920 ;
        RECT 10.270 0.740 10.400 0.920 ;
        RECT 11.230 0.560 11.360 0.920 ;
        RECT 13.150 0.560 13.280 0.920 ;
        RECT 2.505 0.260 2.805 0.560 ;
        RECT 5.385 0.260 5.685 0.560 ;
        RECT 8.265 0.260 8.565 0.560 ;
        RECT 11.145 0.260 11.445 0.560 ;
        RECT 13.065 0.260 13.365 0.560 ;
      LAYER Metal1 ;
        RECT 2.575 5.630 8.545 5.790 ;
        RECT 8.815 5.630 11.425 5.790 ;
        RECT 2.575 4.790 2.735 5.630 ;
        RECT 8.815 5.130 8.975 5.630 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 2.045 4.630 2.785 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 4.975 4.330 5.135 4.630 ;
        RECT 7.855 4.330 8.015 4.630 ;
        RECT 4.925 4.170 5.185 4.330 ;
        RECT 6.365 4.170 8.015 4.330 ;
        RECT 0.175 3.490 8.545 3.650 ;
        RECT 0.175 1.150 0.335 3.490 ;
        RECT 4.925 2.530 7.585 2.690 ;
        RECT 1.565 2.050 3.745 2.210 ;
        RECT 4.975 1.150 5.135 2.530 ;
        RECT 6.365 1.390 8.015 1.550 ;
        RECT 7.855 1.150 8.015 1.390 ;
        RECT 8.815 1.150 8.975 4.630 ;
        RECT 11.695 1.550 11.855 4.630 ;
        RECT 10.205 1.390 12.335 1.550 ;
        RECT 11.695 1.150 11.855 1.390 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 8.765 0.990 11.375 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 11.215 0.490 11.375 0.990 ;
        RECT 12.175 0.490 12.335 1.390 ;
        RECT 2.095 0.330 8.545 0.490 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 12.175 0.330 13.345 0.490 ;
  END
END DFQD1_2

#--------EOF---------

MACRO DFQD1_3
  CLASS CORE ;
  FOREIGN DFQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.142350 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.510 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.325 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 1.615 2.210 1.775 3.490 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 1.150 12.815 4.630 ;
        RECT 12.605 0.990 12.865 1.150 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 10.735 0.150 10.895 0.990 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 3.055 4.790 3.215 5.970 ;
        RECT 10.735 5.130 10.895 5.970 ;
        RECT 10.685 4.970 10.945 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 13.150 5.200 13.280 5.380 ;
        RECT 5.470 4.400 5.600 4.925 ;
        RECT 0.670 3.155 0.800 4.100 ;
        RECT 3.550 3.240 3.680 4.390 ;
        RECT 5.385 4.100 5.685 4.400 ;
        RECT 6.430 3.720 6.560 4.925 ;
        RECT 7.390 4.400 7.520 4.510 ;
        RECT 7.305 4.100 7.605 4.400 ;
        RECT 6.345 3.420 6.645 3.720 ;
        RECT 2.025 3.155 2.325 3.240 ;
        RECT 0.670 3.025 2.325 3.155 ;
        RECT 0.670 1.620 0.800 3.025 ;
        RECT 2.025 2.940 2.325 3.025 ;
        RECT 3.465 2.940 3.765 3.240 ;
        RECT 5.385 2.940 5.685 3.240 ;
        RECT 1.065 2.675 1.365 2.760 ;
        RECT 3.550 2.675 3.680 2.940 ;
        RECT 1.065 2.545 3.680 2.675 ;
        RECT 1.065 2.460 1.365 2.545 ;
        RECT 3.550 1.325 3.680 1.505 ;
        RECT 5.470 1.165 5.600 2.940 ;
        RECT 6.430 1.620 6.560 3.420 ;
        RECT 7.390 2.760 7.520 4.100 ;
        RECT 7.785 2.940 8.085 3.240 ;
        RECT 7.305 2.460 7.605 2.760 ;
        RECT 6.345 1.320 6.645 1.620 ;
        RECT 7.390 1.375 7.520 2.460 ;
        RECT 7.870 2.195 8.000 2.940 ;
        RECT 8.350 2.760 8.480 4.225 ;
        RECT 9.310 3.240 9.440 4.925 ;
        RECT 9.225 2.940 9.525 3.240 ;
        RECT 8.265 2.460 8.565 2.760 ;
        RECT 7.870 2.065 8.480 2.195 ;
        RECT 6.430 1.165 6.560 1.320 ;
        RECT 8.350 1.295 8.480 2.065 ;
        RECT 9.310 1.165 9.440 1.345 ;
        RECT 10.270 1.165 10.400 4.925 ;
        RECT 11.230 2.280 11.360 4.100 ;
        RECT 11.145 1.980 11.445 2.280 ;
        RECT 11.230 1.620 11.360 1.980 ;
        RECT 13.150 1.620 13.280 4.100 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 7.390 0.740 7.520 0.920 ;
        RECT 8.350 0.740 8.480 0.920 ;
        RECT 9.310 0.560 9.440 0.920 ;
        RECT 3.465 0.260 3.765 0.560 ;
        RECT 9.225 0.260 9.525 0.560 ;
        RECT 10.270 0.475 10.400 0.920 ;
        RECT 11.230 0.740 11.360 0.920 ;
        RECT 11.625 0.475 11.925 0.560 ;
        RECT 13.150 0.475 13.280 0.920 ;
        RECT 10.270 0.345 13.280 0.475 ;
        RECT 11.625 0.260 11.925 0.345 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 4.925 4.630 7.535 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 8.765 4.630 11.375 4.790 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 0.175 2.690 0.335 4.630 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 7.375 4.330 7.535 4.630 ;
        RECT 2.095 4.170 5.665 4.330 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 2.095 3.170 2.255 4.170 ;
        RECT 7.855 3.650 8.015 4.630 ;
        RECT 6.365 3.490 8.015 3.650 ;
        RECT 2.045 3.010 2.305 3.170 ;
        RECT 3.485 3.010 9.505 3.170 ;
        RECT 0.175 2.530 1.345 2.690 ;
        RECT 0.175 1.150 0.335 2.530 ;
        RECT 2.095 1.150 2.255 3.010 ;
        RECT 4.975 2.530 7.585 2.690 ;
        RECT 8.285 2.530 8.545 2.690 ;
        RECT 4.975 1.150 5.135 2.530 ;
        RECT 6.365 1.390 8.015 1.550 ;
        RECT 7.855 1.150 8.015 1.390 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 8.335 0.490 8.495 2.530 ;
        RECT 11.215 2.210 11.375 4.630 ;
        RECT 8.815 2.050 11.425 2.210 ;
        RECT 8.815 1.150 8.975 2.050 ;
        RECT 11.695 1.150 11.855 4.630 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 11.695 0.490 11.855 0.990 ;
        RECT 2.095 0.330 9.505 0.490 ;
        RECT 11.645 0.330 11.905 0.490 ;
  END
END DFQD1_3

#--------EOF---------

MACRO FILL1
  CLASS CORE ;
  FOREIGN FILL1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.340 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.340 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 0.340 6.270 ;
    END
  END vdd
END FILL1

#--------EOF---------

MACRO FILL2
  CLASS CORE ;
  FOREIGN FILL2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.680 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.680 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 0.680 6.270 ;
    END
  END vdd
END FILL2

#--------EOF---------

MACRO FILL4
  CLASS CORE ;
  FOREIGN FILL4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.360 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 1.360 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.360 6.270 ;
    END
  END vdd
END FILL4

#--------EOF---------

MACRO FILL8
  CLASS CORE ;
  FOREIGN FILL8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END FILL8

#--------EOF---------

MACRO INVD1
  CLASS CORE ;
  FOREIGN INVD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
END INVD1

#--------EOF---------

MACRO INVD1_1
  CLASS CORE ;
  FOREIGN INVD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
END INVD1_1

#--------EOF---------

MACRO INVD1_2
  CLASS CORE ;
  FOREIGN INVD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
END INVD1_2

#--------EOF---------

MACRO INVD1_3
  CLASS CORE ;
  FOREIGN INVD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
END INVD1_3

#--------EOF---------

MACRO MUX2D1
  CLASS CORE ;
  FOREIGN MUX2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.645 5.600 5.775 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 3.550 4.470 3.680 4.650 ;
        RECT 5.470 4.400 5.600 4.650 ;
        RECT 5.385 4.100 5.685 4.400 ;
        RECT 5.385 1.980 5.685 2.280 ;
        RECT 4.425 1.535 4.725 1.620 ;
        RECT 5.470 1.535 5.600 1.980 ;
        RECT 0.670 1.270 0.800 1.450 ;
        RECT 4.425 1.405 5.600 1.535 ;
        RECT 4.425 1.320 4.725 1.405 ;
        RECT 5.470 1.270 5.600 1.405 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 5.455 2.210 5.615 4.170 ;
        RECT 5.405 2.050 5.665 2.210 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 4.495 0.490 4.655 1.390 ;
        RECT 0.605 0.330 4.655 0.490 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.050 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.183950 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 3.635 2.720 4.290 ;
        RECT 2.110 3.505 2.720 3.635 ;
        RECT 2.110 2.195 2.240 3.505 ;
        RECT 2.505 2.195 2.805 2.280 ;
        RECT 2.110 2.065 2.805 2.195 ;
        RECT 2.505 1.980 2.805 2.065 ;
        RECT 2.590 1.425 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 1.390 2.735 2.050 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830550 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 1.150 7.055 4.630 ;
        RECT 6.845 0.990 7.105 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 2.045 4.630 2.305 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.985 5.775 3.285 5.860 ;
        RECT 0.670 5.645 3.285 5.775 ;
        RECT 0.670 5.200 0.800 5.645 ;
        RECT 2.985 5.560 3.285 5.645 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 4.470 0.800 4.650 ;
        RECT 1.065 3.420 1.365 3.720 ;
        RECT 3.945 3.635 4.245 3.720 ;
        RECT 6.430 3.635 6.560 4.430 ;
        RECT 3.945 3.505 6.560 3.635 ;
        RECT 3.945 3.420 4.245 3.505 ;
        RECT 1.150 2.280 1.280 3.420 ;
        RECT 2.505 2.675 2.805 2.760 ;
        RECT 3.945 2.675 4.245 2.760 ;
        RECT 2.505 2.545 6.560 2.675 ;
        RECT 2.505 2.460 2.805 2.545 ;
        RECT 3.945 2.460 4.245 2.545 ;
        RECT 1.065 1.980 1.365 2.280 ;
        RECT 6.430 1.620 6.560 2.545 ;
        RECT 3.550 1.270 3.680 1.450 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 4.905 0.475 5.205 0.560 ;
        RECT 3.550 0.345 5.205 0.475 ;
        RECT 4.905 0.260 5.205 0.345 ;
      LAYER Metal1 ;
        RECT 3.005 5.630 5.135 5.790 ;
        RECT 4.975 5.130 5.135 5.630 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.175 2.690 0.335 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 3.650 1.295 4.630 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 0.175 2.530 2.785 2.690 ;
        RECT 0.175 1.150 0.335 2.530 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 1.135 1.150 1.295 2.050 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 4.015 3.650 4.175 4.970 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 4.015 2.690 4.175 3.490 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 4.015 1.150 4.175 2.530 ;
        RECT 4.975 1.150 5.135 4.970 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 4.925 0.330 5.185 0.490 ;
  END
END MUX2D1

#--------EOF---------

MACRO MUX2D1_1
  CLASS CORE ;
  FOREIGN MUX2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 3.155 2.720 4.650 ;
        RECT 4.510 3.240 4.640 4.650 ;
        RECT 2.985 3.155 3.285 3.240 ;
        RECT 1.630 3.025 3.285 3.155 ;
        RECT 1.630 1.270 1.760 3.025 ;
        RECT 2.985 2.940 3.285 3.025 ;
        RECT 4.425 2.940 4.725 3.240 ;
        RECT 4.510 1.270 4.640 2.940 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 3.010 4.705 3.170 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.183950 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.290 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.425 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830550 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.545 5.560 1.845 5.860 ;
        RECT 1.630 5.200 1.760 5.560 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 3.720 1.760 4.650 ;
        RECT 4.905 4.315 5.205 4.400 ;
        RECT 6.430 4.315 6.560 4.430 ;
        RECT 4.905 4.185 6.560 4.315 ;
        RECT 4.905 4.100 5.205 4.185 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.270 2.720 1.980 ;
        RECT 6.430 1.620 6.560 4.185 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 6.430 0.560 6.560 0.920 ;
        RECT 6.345 0.260 6.645 0.560 ;
      LAYER Metal1 ;
        RECT 1.565 5.630 5.135 5.790 ;
        RECT 4.975 5.130 5.135 5.630 ;
        RECT 2.045 4.970 4.655 5.130 ;
        RECT 4.925 4.970 5.615 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.575 4.630 3.265 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 1.615 2.210 1.775 3.490 ;
        RECT 2.575 2.690 2.735 4.630 ;
        RECT 4.495 4.330 4.655 4.970 ;
        RECT 4.495 4.170 5.185 4.330 ;
        RECT 2.575 2.530 3.215 2.690 ;
        RECT 1.615 2.050 2.785 2.210 ;
        RECT 3.055 1.150 3.215 2.530 ;
        RECT 5.455 1.150 5.615 4.970 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.615 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 2.095 0.330 6.625 0.490 ;
  END
END MUX2D1_1

#--------EOF---------

MACRO MUX2D1_2
  CLASS CORE ;
  FOREIGN MUX2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.645 5.600 5.775 ;
        RECT 0.670 5.200 0.800 5.645 ;
        RECT 5.470 5.200 5.600 5.645 ;
        RECT 0.670 4.470 0.800 4.650 ;
        RECT 4.425 2.195 4.725 2.280 ;
        RECT 5.470 2.195 5.600 4.650 ;
        RECT 3.550 2.065 5.600 2.195 ;
        RECT 3.550 1.270 3.680 2.065 ;
        RECT 4.425 1.980 4.725 2.065 ;
        RECT 5.470 1.270 5.600 2.065 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.183950 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.290 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.425 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830550 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 1.150 7.055 4.630 ;
        RECT 6.845 0.990 7.105 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 5.935 0.150 6.095 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 2.045 4.630 2.305 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.065 3.420 1.365 3.720 ;
        RECT 2.985 3.420 3.285 3.720 ;
        RECT 1.150 2.280 1.280 3.420 ;
        RECT 3.070 2.280 3.200 3.420 ;
        RECT 3.550 2.760 3.680 4.650 ;
        RECT 3.465 2.460 3.765 2.760 ;
        RECT 1.065 1.980 1.365 2.280 ;
        RECT 2.985 1.980 3.285 2.280 ;
        RECT 6.430 1.620 6.560 4.430 ;
        RECT 0.670 1.270 0.800 1.450 ;
        RECT 4.425 0.920 4.725 1.220 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.465 0.475 3.765 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 0.670 0.345 4.640 0.475 ;
        RECT 4.905 0.475 5.205 0.560 ;
        RECT 6.430 0.475 6.560 0.920 ;
        RECT 4.905 0.345 6.560 0.475 ;
        RECT 3.465 0.260 3.765 0.345 ;
        RECT 4.905 0.260 5.205 0.345 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.815 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.655 3.170 0.815 4.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 3.650 1.295 4.630 ;
        RECT 3.055 3.650 3.215 4.630 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 4.015 3.170 4.175 4.970 ;
        RECT 0.175 3.010 4.175 3.170 ;
        RECT 0.175 1.150 0.335 3.010 ;
        RECT 3.485 2.530 3.745 2.690 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 1.135 1.150 1.295 2.050 ;
        RECT 3.055 1.150 3.215 2.050 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.535 0.490 3.695 2.530 ;
        RECT 4.015 1.150 4.175 3.010 ;
        RECT 4.975 1.150 5.135 4.970 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.445 0.990 5.185 1.150 ;
        RECT 4.015 0.490 4.175 0.990 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 4.015 0.330 5.185 0.490 ;
  END
END MUX2D1_2

#--------EOF---------

MACRO MUX2D1_3
  CLASS CORE ;
  FOREIGN MUX2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.645 4.640 5.775 ;
        RECT 1.630 5.200 1.760 5.645 ;
        RECT 4.510 5.200 4.640 5.645 ;
        RECT 1.630 4.470 1.760 4.650 ;
        RECT 4.510 3.635 4.640 4.650 ;
        RECT 4.030 3.505 4.640 3.635 ;
        RECT 4.030 2.195 4.160 3.505 ;
        RECT 4.030 2.065 4.640 2.195 ;
        RECT 2.590 1.270 2.720 1.450 ;
        RECT 4.510 1.270 4.640 2.065 ;
        RECT 2.590 0.560 2.720 0.920 ;
        RECT 2.505 0.475 2.805 0.560 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 2.505 0.345 4.640 0.475 ;
        RECT 2.505 0.260 2.805 0.345 ;
      LAYER Metal1 ;
        RECT 2.575 0.490 2.735 1.150 ;
        RECT 2.525 0.330 2.785 0.490 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.183950 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.290 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.425 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830550 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 2.590 4.400 2.720 4.650 ;
        RECT 2.505 4.100 2.805 4.400 ;
        RECT 2.590 3.635 2.720 4.100 ;
        RECT 1.630 3.505 2.720 3.635 ;
        RECT 1.630 1.270 1.760 3.505 ;
        RECT 2.985 3.420 3.285 3.720 ;
        RECT 3.070 2.280 3.200 3.420 ;
        RECT 4.425 3.155 4.725 3.240 ;
        RECT 6.430 3.155 6.560 4.430 ;
        RECT 4.425 3.025 6.560 3.155 ;
        RECT 4.425 2.940 4.725 3.025 ;
        RECT 2.985 1.980 3.285 2.280 ;
        RECT 6.430 1.620 6.560 3.025 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.575 4.970 3.695 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 2.095 3.170 2.255 4.970 ;
        RECT 2.575 4.330 2.735 4.970 ;
        RECT 3.535 4.790 3.695 4.970 ;
        RECT 4.975 4.790 5.135 4.970 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.535 4.630 5.135 4.790 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 3.055 3.650 3.215 4.630 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 2.095 3.010 4.705 3.170 ;
        RECT 2.095 1.150 2.255 3.010 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.055 1.150 3.215 2.050 ;
        RECT 4.975 1.150 5.135 4.630 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
  END
END MUX2D1_3

#--------EOF---------

MACRO ND2D1
  CLASS CORE ;
  FOREIGN ND2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.308500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 2.255 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
    END
  END vdd
END ND2D1

#--------EOF---------

MACRO ND2D1_1
  CLASS CORE ;
  FOREIGN ND2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.308500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 4.630 1.345 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 2.045 4.630 2.305 4.790 ;
    END
  END vdd
END ND2D1_1

#--------EOF---------

MACRO ND2D1_2
  CLASS CORE ;
  FOREIGN ND2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END ND2D1_2

#--------EOF---------

MACRO ND2D1_3
  CLASS CORE ;
  FOREIGN ND2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 2.305 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END ND2D1_3

#--------EOF---------

MACRO ND3D1
  CLASS CORE ;
  FOREIGN ND3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.930000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 4.630 3.265 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 1.150 2.255 4.170 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 0.175 0.330 3.215 0.490 ;
  END
END ND3D1

#--------EOF---------

MACRO ND3D1_1
  CLASS CORE ;
  FOREIGN ND3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.930000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.400 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.400 6.270 ;
    END
  END vdd
END ND3D1_1

#--------EOF---------

MACRO ND3D1_2
  CLASS CORE ;
  FOREIGN ND3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.760 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.930000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 4.015 0.490 4.175 0.990 ;
        RECT 0.175 0.330 4.175 0.490 ;
  END
END ND3D1_2

#--------EOF---------

MACRO ND3D1_3
  CLASS CORE ;
  FOREIGN ND3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.260000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 3.265 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 0.175 0.330 3.215 0.490 ;
  END
END ND3D1_3

#--------EOF---------

MACRO ND4D1
  CLASS CORE ;
  FOREIGN ND4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.100 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.620 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.551500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 3.055 1.150 3.215 4.170 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 4.015 0.490 4.175 0.990 ;
        RECT 0.175 0.330 4.175 0.490 ;
  END
END ND4D1

#--------EOF---------

MACRO ND4D1_1
  CLASS CORE ;
  FOREIGN ND4D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.551500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 4.225 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 4.015 1.150 4.175 4.170 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.100 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.620 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 4.975 4.790 5.135 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 0.175 0.330 5.135 0.490 ;
  END
END ND4D1_1

#--------EOF---------

MACRO ND4D1_2
  CLASS CORE ;
  FOREIGN ND4D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.221500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 3.265 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.135 0.990 4.225 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
END ND4D1_2

#--------EOF---------

MACRO ND4D1_3
  CLASS CORE ;
  FOREIGN ND4D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.221500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 1.135 4.170 5.135 4.330 ;
        RECT 4.975 1.150 5.135 4.170 ;
        RECT 4.925 0.990 5.185 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.100 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.620 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 3.055 4.790 3.215 5.970 ;
        RECT 4.975 4.790 5.135 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 3.265 1.150 ;
  END
END ND4D1_3

#--------EOF---------

MACRO NR2D1
  CLASS CORE ;
  FOREIGN NR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.202500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 1.295 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 2.095 4.790 2.255 5.970 ;
        RECT 2.045 4.630 2.305 4.790 ;
    END
  END vdd
END NR2D1

#--------EOF---------

MACRO NR2D1_1
  CLASS CORE ;
  FOREIGN NR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.202500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 4.630 2.305 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
    END
  END vdd
END NR2D1_1

#--------EOF---------

MACRO NR2D1_2
  CLASS CORE ;
  FOREIGN NR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.412500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END NR2D1_2

#--------EOF---------

MACRO NR2D1_3
  CLASS CORE ;
  FOREIGN NR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.412500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 0.125 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END
  END vdd
END NR2D1_3

#--------EOF---------

MACRO NR3D1
  CLASS CORE ;
  FOREIGN NR3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.889500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 3.265 1.150 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 4.510 3.155 4.640 4.100 ;
        RECT 6.430 3.635 6.560 4.100 ;
        RECT 5.470 3.505 6.560 3.635 ;
        RECT 5.470 3.155 5.600 3.505 ;
        RECT 4.510 3.025 5.600 3.155 ;
        RECT 1.545 2.195 1.845 2.280 ;
        RECT 4.510 2.195 4.640 3.025 ;
        RECT 0.670 2.065 4.640 2.195 ;
        RECT 0.670 1.620 0.800 2.065 ;
        RECT 1.545 1.980 1.845 2.065 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 2.590 3.720 2.720 4.100 ;
        RECT 2.505 3.420 2.805 3.720 ;
        RECT 6.825 3.635 7.125 3.720 ;
        RECT 8.350 3.635 8.480 4.100 ;
        RECT 6.825 3.505 8.480 3.635 ;
        RECT 6.825 3.420 7.125 3.505 ;
        RECT 6.910 2.675 7.040 3.420 ;
        RECT 5.950 2.545 7.040 2.675 ;
        RECT 2.590 1.620 2.720 1.800 ;
        RECT 5.950 1.535 6.080 2.545 ;
        RECT 4.990 1.405 6.080 1.535 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 4.990 0.475 5.120 1.405 ;
        RECT 2.590 0.345 5.120 0.475 ;
      LAYER Metal1 ;
        RECT 2.525 3.490 7.105 3.650 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.635 0.885 3.720 ;
        RECT 1.630 3.635 1.760 4.100 ;
        RECT 0.585 3.505 1.760 3.635 ;
        RECT 0.585 3.420 0.885 3.505 ;
        RECT 1.630 1.620 1.760 1.800 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 0.585 0.345 1.760 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
      LAYER Metal1 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 0.490 0.815 3.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 1.615 4.790 1.775 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.630 8.065 4.790 ;
        RECT 8.335 4.630 9.025 4.790 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 3.055 4.170 4.175 4.330 ;
        RECT 5.935 4.330 6.095 4.630 ;
        RECT 8.335 4.330 8.495 4.630 ;
        RECT 5.935 4.170 8.495 4.330 ;
  END
END NR3D1

#--------EOF---------

MACRO NR3D1_1
  CLASS CORE ;
  FOREIGN NR3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.540 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.889500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.550 1.295 4.630 ;
        RECT 1.135 1.390 3.215 1.550 ;
        RECT 1.135 1.150 1.295 1.390 ;
        RECT 3.055 1.150 3.215 1.390 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 1.545 2.195 1.845 2.280 ;
        RECT 5.470 2.195 5.600 4.100 ;
        RECT 7.390 2.195 7.520 4.100 ;
        RECT 1.545 2.065 7.520 2.195 ;
        RECT 1.545 1.980 1.845 2.065 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 3.550 3.720 3.680 4.100 ;
        RECT 3.465 3.420 3.765 3.720 ;
        RECT 3.550 1.620 3.680 1.800 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 3.465 0.475 3.765 0.560 ;
        RECT 9.310 0.475 9.440 4.100 ;
        RECT 3.465 0.345 9.440 0.475 ;
        RECT 3.465 0.260 3.765 0.345 ;
      LAYER Metal1 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 3.535 0.490 3.695 3.490 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 3.635 0.800 4.100 ;
        RECT 1.630 3.635 1.760 4.100 ;
        RECT 0.670 3.505 1.760 3.635 ;
        RECT 0.670 2.280 0.800 3.505 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 10.540 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 10.540 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.330 1.775 4.970 ;
        RECT 2.095 4.970 8.975 5.130 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 8.815 4.790 8.975 4.970 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.965 4.630 5.185 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 1.615 4.170 3.215 4.330 ;
        RECT 6.895 4.330 7.055 4.630 ;
        RECT 9.775 4.330 9.935 4.630 ;
        RECT 6.895 4.170 9.935 4.330 ;
  END
END NR3D1_1

#--------EOF---------

MACRO NR3D1_2
  CLASS CORE ;
  FOREIGN NR3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.889500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 0.125 0.990 2.305 1.150 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 4.510 3.155 4.640 4.100 ;
        RECT 6.430 3.635 6.560 4.100 ;
        RECT 5.470 3.505 6.560 3.635 ;
        RECT 5.470 3.155 5.600 3.505 ;
        RECT 4.510 3.025 5.600 3.155 ;
        RECT 0.585 2.195 0.885 2.280 ;
        RECT 4.510 2.195 4.640 3.025 ;
        RECT 0.585 2.065 4.640 2.195 ;
        RECT 0.585 1.980 0.885 2.065 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 2.590 3.720 2.720 4.100 ;
        RECT 2.505 3.420 2.805 3.720 ;
        RECT 8.350 2.760 8.480 4.100 ;
        RECT 8.265 2.460 8.565 2.760 ;
        RECT 2.590 1.620 2.720 1.800 ;
        RECT 2.590 0.560 2.720 0.920 ;
        RECT 2.505 0.260 2.805 0.560 ;
      LAYER Metal1 ;
        RECT 2.525 3.490 2.785 3.650 ;
        RECT 2.575 0.490 2.735 3.490 ;
        RECT 5.935 2.530 8.545 2.690 ;
        RECT 5.935 1.550 6.095 2.530 ;
        RECT 4.975 1.390 6.095 1.550 ;
        RECT 4.975 0.490 5.135 1.390 ;
        RECT 2.525 0.330 5.135 0.490 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.143000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 3.720 1.760 4.100 ;
        RECT 1.545 3.420 1.845 3.720 ;
      LAYER Metal1 ;
        RECT 1.615 3.650 1.775 4.330 ;
        RECT 1.565 3.490 1.825 3.650 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.920 0.800 4.100 ;
        RECT 1.630 1.620 1.760 1.800 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 1.615 4.790 1.775 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.630 8.065 4.790 ;
        RECT 8.335 4.630 9.025 4.790 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 3.055 4.170 4.175 4.330 ;
        RECT 5.935 4.330 6.095 4.630 ;
        RECT 8.335 4.330 8.495 4.630 ;
        RECT 5.935 4.170 8.495 4.330 ;
  END
END NR3D1_2

#--------EOF---------

MACRO NR3D1_3
  CLASS CORE ;
  FOREIGN NR3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.889500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.735 4.790 ;
        RECT 2.575 1.550 2.735 4.630 ;
        RECT 1.135 1.390 2.735 1.550 ;
        RECT 1.135 1.150 1.295 1.390 ;
        RECT 2.575 1.150 2.735 1.390 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.575 0.990 3.265 1.150 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 2.985 2.195 3.285 2.280 ;
        RECT 4.510 2.195 4.640 4.100 ;
        RECT 6.430 2.195 6.560 4.100 ;
        RECT 2.590 2.065 6.560 2.195 ;
        RECT 2.590 1.620 2.720 2.065 ;
        RECT 2.985 1.980 3.285 2.065 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 3.055 2.210 3.215 2.690 ;
        RECT 3.005 2.050 3.265 2.210 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 0.670 1.620 0.800 4.100 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 8.350 0.475 8.480 4.100 ;
        RECT 0.585 0.345 8.480 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
      LAYER Metal1 ;
        RECT 0.655 0.490 0.815 1.150 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.377000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 1.630 3.635 1.760 4.100 ;
        RECT 2.590 3.635 2.720 4.100 ;
        RECT 1.630 3.505 2.720 3.635 ;
        RECT 1.630 2.280 1.760 3.505 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.150 2.255 0.990 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.175 4.970 4.175 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 4.015 4.790 4.175 4.970 ;
        RECT 5.935 4.970 8.975 5.130 ;
        RECT 5.935 4.790 6.095 4.970 ;
        RECT 8.815 4.790 8.975 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 7.855 4.330 8.015 4.630 ;
        RECT 3.055 4.170 8.015 4.330 ;
  END
END NR3D1_3

#--------EOF---------

MACRO NR4D1
  CLASS CORE ;
  FOREIGN NR4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.260 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.668300 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 4.225 1.150 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 8.350 3.155 8.480 4.100 ;
        RECT 10.270 3.635 10.400 4.100 ;
        RECT 9.310 3.505 10.400 3.635 ;
        RECT 9.310 3.155 9.440 3.505 ;
        RECT 8.350 3.025 9.440 3.155 ;
        RECT 4.425 2.195 4.725 2.280 ;
        RECT 8.350 2.195 8.480 3.025 ;
        RECT 4.425 2.065 8.480 2.195 ;
        RECT 4.425 1.980 4.725 2.065 ;
        RECT 4.510 1.375 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 4.510 2.675 4.640 4.100 ;
        RECT 12.190 3.720 12.320 4.100 ;
        RECT 7.785 3.420 8.085 3.720 ;
        RECT 12.105 3.420 12.405 3.720 ;
        RECT 7.870 2.675 8.000 3.420 ;
        RECT 4.030 2.545 8.000 2.675 ;
        RECT 4.030 2.195 4.160 2.545 ;
        RECT 3.550 2.065 4.160 2.195 ;
        RECT 3.550 1.375 3.680 2.065 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 7.805 3.490 12.385 3.650 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 6.430 3.720 6.560 4.100 ;
        RECT 3.945 3.635 4.245 3.720 ;
        RECT 2.590 3.505 4.245 3.635 ;
        RECT 2.590 3.155 2.720 3.505 ;
        RECT 3.945 3.420 4.245 3.505 ;
        RECT 6.345 3.420 6.645 3.720 ;
        RECT 1.630 3.025 2.720 3.155 ;
        RECT 1.630 2.195 1.760 3.025 ;
        RECT 0.670 2.065 1.760 2.195 ;
        RECT 0.670 1.375 0.800 2.065 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 3.965 3.490 6.625 3.650 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.635 0.885 3.720 ;
        RECT 1.630 3.635 1.760 4.100 ;
        RECT 0.585 3.505 1.760 3.635 ;
        RECT 0.585 3.420 0.885 3.505 ;
        RECT 1.630 1.375 1.760 1.555 ;
        RECT 0.585 0.475 0.885 0.560 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 0.585 0.345 1.760 0.475 ;
        RECT 0.585 0.260 0.885 0.345 ;
      LAYER Metal1 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 0.490 0.815 3.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 7.305 4.900 7.605 5.200 ;
        RECT 7.390 4.400 7.520 4.900 ;
        RECT 7.305 4.100 7.605 4.400 ;
      LAYER Metal1 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 7.325 4.970 9.935 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 1.615 4.790 1.775 4.970 ;
        RECT 9.775 4.790 9.935 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.630 3.265 4.790 ;
        RECT 4.925 4.630 6.575 4.790 ;
        RECT 6.845 4.630 11.905 4.790 ;
        RECT 12.175 4.630 12.865 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 5.935 4.330 6.095 4.630 ;
        RECT 2.095 4.170 6.095 4.330 ;
        RECT 6.415 4.330 6.575 4.630 ;
        RECT 7.855 4.330 8.015 4.630 ;
        RECT 12.175 4.330 12.335 4.630 ;
        RECT 6.415 4.170 7.585 4.330 ;
        RECT 7.855 4.170 12.335 4.330 ;
  END
END NR4D1

#--------EOF---------

MACRO NR4D1_1
  CLASS CORE ;
  FOREIGN NR4D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.668300 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 1.085 0.990 3.265 1.150 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 7.390 5.200 7.520 5.380 ;
        RECT 9.310 5.200 9.440 5.380 ;
        RECT 7.390 3.155 7.520 4.100 ;
        RECT 9.310 3.635 9.440 4.100 ;
        RECT 8.350 3.505 9.440 3.635 ;
        RECT 8.350 3.155 8.480 3.505 ;
        RECT 7.390 3.025 8.480 3.155 ;
        RECT 3.465 2.195 3.765 2.280 ;
        RECT 7.390 2.195 7.520 3.025 ;
        RECT 3.465 2.065 7.520 2.195 ;
        RECT 3.465 1.980 3.765 2.065 ;
        RECT 3.550 1.375 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 11.230 5.200 11.360 5.380 ;
        RECT 3.550 2.675 3.680 4.100 ;
        RECT 11.230 3.720 11.360 4.100 ;
        RECT 6.825 3.420 7.125 3.720 ;
        RECT 11.145 3.420 11.445 3.720 ;
        RECT 6.910 2.675 7.040 3.420 ;
        RECT 3.070 2.545 7.040 2.675 ;
        RECT 3.070 2.195 3.200 2.545 ;
        RECT 2.590 2.065 3.200 2.195 ;
        RECT 2.590 1.375 2.720 2.065 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 6.845 3.490 11.425 3.650 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 2.590 3.635 2.720 4.100 ;
        RECT 5.470 3.720 5.600 4.100 ;
        RECT 2.985 3.635 3.285 3.720 ;
        RECT 1.630 3.505 3.285 3.635 ;
        RECT 1.630 1.375 1.760 3.505 ;
        RECT 2.985 3.420 3.285 3.505 ;
        RECT 5.385 3.420 5.685 3.720 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 3.005 3.490 5.665 3.650 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.645 1.760 5.775 ;
        RECT 0.670 5.200 0.800 5.645 ;
        RECT 1.630 5.200 1.760 5.645 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 1.630 3.920 1.760 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.375 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 6.345 4.900 6.645 5.200 ;
        RECT 6.430 4.400 6.560 4.900 ;
        RECT 6.345 4.100 6.645 4.400 ;
      LAYER Metal1 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 6.365 4.970 8.975 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.330 1.775 4.970 ;
        RECT 8.815 4.790 8.975 4.970 ;
        RECT 3.965 4.630 5.615 4.790 ;
        RECT 5.885 4.630 10.945 4.790 ;
        RECT 11.215 4.630 11.905 4.790 ;
        RECT 4.975 4.330 5.135 4.630 ;
        RECT 1.615 4.170 5.135 4.330 ;
        RECT 5.455 4.330 5.615 4.630 ;
        RECT 6.895 4.330 7.055 4.630 ;
        RECT 11.215 4.330 11.375 4.630 ;
        RECT 5.455 4.170 6.625 4.330 ;
        RECT 6.895 4.170 11.375 4.330 ;
  END
END NR4D1_1

#--------EOF---------

MACRO NR4D1_2
  CLASS CORE ;
  FOREIGN NR4D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.260 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.668300 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 1.150 4.175 4.630 ;
        RECT 1.085 0.990 4.225 1.150 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 8.350 5.200 8.480 5.380 ;
        RECT 10.270 5.200 10.400 5.380 ;
        RECT 8.350 3.155 8.480 4.100 ;
        RECT 10.270 3.635 10.400 4.100 ;
        RECT 9.310 3.505 10.400 3.635 ;
        RECT 9.310 3.155 9.440 3.505 ;
        RECT 8.350 3.025 9.440 3.155 ;
        RECT 1.545 2.195 1.845 2.280 ;
        RECT 8.350 2.195 8.480 3.025 ;
        RECT 1.545 2.065 8.480 2.195 ;
        RECT 1.545 1.980 1.845 2.065 ;
        RECT 1.630 1.375 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 12.190 5.200 12.320 5.380 ;
        RECT 1.630 2.675 1.760 4.100 ;
        RECT 12.190 3.720 12.320 4.100 ;
        RECT 7.785 3.420 8.085 3.720 ;
        RECT 12.105 3.420 12.405 3.720 ;
        RECT 7.870 2.675 8.000 3.420 ;
        RECT 1.150 2.545 8.000 2.675 ;
        RECT 1.150 2.195 1.280 2.545 ;
        RECT 0.670 2.065 1.280 2.195 ;
        RECT 0.670 1.375 0.800 2.065 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 7.805 3.490 12.385 3.650 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 3.465 3.635 3.765 3.720 ;
        RECT 6.430 3.635 6.560 4.100 ;
        RECT 3.465 3.505 6.560 3.635 ;
        RECT 3.465 3.420 3.765 3.505 ;
        RECT 3.550 1.375 3.680 1.555 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 3.465 0.260 3.765 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 3.490 3.745 3.650 ;
        RECT 0.655 0.490 0.815 3.490 ;
        RECT 0.655 0.330 3.745 0.490 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.345150 ;
    PORT
      LAYER GatPoly ;
        RECT 3.465 5.560 3.765 5.860 ;
        RECT 4.425 5.560 4.725 5.860 ;
        RECT 3.550 5.200 3.680 5.560 ;
        RECT 4.510 5.200 4.640 5.560 ;
        RECT 3.550 3.920 3.680 4.100 ;
        RECT 4.510 3.920 4.640 4.100 ;
        RECT 4.510 1.375 4.640 1.555 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.260 4.725 0.560 ;
      LAYER Metal1 ;
        RECT 3.485 5.630 4.705 5.790 ;
        RECT 4.495 0.490 4.655 5.630 ;
        RECT 4.445 0.330 4.705 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 7.305 4.900 7.605 5.200 ;
        RECT 2.505 4.100 2.805 4.400 ;
        RECT 2.590 3.155 2.720 4.100 ;
        RECT 7.390 3.155 7.520 4.900 ;
        RECT 2.590 3.025 7.520 3.155 ;
      LAYER Metal1 ;
        RECT 7.325 4.970 9.935 5.130 ;
        RECT 9.775 4.790 9.935 4.970 ;
        RECT 0.125 4.630 3.265 4.790 ;
        RECT 4.925 4.630 6.145 4.790 ;
        RECT 6.845 4.630 11.905 4.790 ;
        RECT 12.175 4.630 12.865 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 7.855 4.330 8.015 4.630 ;
        RECT 12.175 4.330 12.335 4.630 ;
        RECT 2.095 4.170 2.785 4.330 ;
        RECT 7.855 4.170 12.335 4.330 ;
  END
END NR4D1_2

#--------EOF---------

MACRO OA21D1
  CLASS CORE ;
  FOREIGN OA21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.100 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.620 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 4.495 2.210 4.655 2.690 ;
        RECT 4.445 2.050 4.705 2.210 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.760 0.800 4.100 ;
        RECT 0.585 2.460 0.885 2.760 ;
        RECT 0.670 1.620 0.800 2.460 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.690 0.815 3.170 ;
        RECT 0.605 2.530 0.865 2.690 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.760 1.760 4.100 ;
        RECT 1.545 2.460 1.845 2.760 ;
        RECT 1.630 1.620 1.760 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.690 1.775 3.170 ;
        RECT 1.565 2.530 1.825 2.690 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 3.465 0.920 3.765 1.220 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 2.590 0.345 3.680 0.475 ;
      LAYER Metal1 ;
        RECT 0.175 4.970 4.175 5.130 ;
        RECT 0.175 4.790 0.335 4.970 ;
        RECT 4.015 4.790 4.175 4.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 0.175 4.170 1.295 4.330 ;
        RECT 0.175 2.210 0.335 4.170 ;
        RECT 0.175 2.050 2.785 2.210 ;
        RECT 0.175 1.150 0.335 2.050 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.485 0.990 4.225 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 1.135 0.330 5.135 0.490 ;
  END
END OA21D1

#--------EOF---------

MACRO OA21D1_1
  CLASS CORE ;
  FOREIGN OA21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.760 2.720 4.100 ;
        RECT 2.505 2.460 2.805 2.760 ;
        RECT 2.590 1.620 2.720 2.460 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.690 2.735 3.170 ;
        RECT 2.525 2.530 2.785 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 1.150 4.175 4.630 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.985 2.195 3.285 2.280 ;
        RECT 4.510 2.195 4.640 4.100 ;
        RECT 2.985 2.065 4.640 2.195 ;
        RECT 2.985 1.980 3.285 2.065 ;
        RECT 4.510 1.620 4.640 2.065 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 2.210 2.255 4.170 ;
        RECT 2.095 2.050 3.265 2.210 ;
        RECT 2.095 1.150 2.255 2.050 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OA21D1_1

#--------EOF---------

MACRO OA21D1_2
  CLASS CORE ;
  FOREIGN OA21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.760 1.760 4.100 ;
        RECT 1.545 2.460 1.845 2.760 ;
        RECT 1.630 1.620 1.760 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.690 1.775 3.170 ;
        RECT 1.565 2.530 1.825 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.760 2.720 4.100 ;
        RECT 2.505 2.460 2.805 2.760 ;
        RECT 2.590 1.620 2.720 2.460 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.690 2.735 3.170 ;
        RECT 2.525 2.530 2.785 2.690 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.465 4.560 3.765 4.860 ;
        RECT 3.550 1.220 3.680 4.560 ;
        RECT 3.465 0.920 3.765 1.220 ;
      LAYER Metal1 ;
        RECT 3.485 4.630 4.225 4.790 ;
        RECT 3.485 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.280 4.640 4.100 ;
        RECT 4.425 1.980 4.725 2.280 ;
        RECT 4.510 1.620 4.640 1.980 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 4.330 0.335 4.630 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 0.175 4.170 3.215 4.330 ;
        RECT 1.135 2.210 1.295 4.170 ;
        RECT 1.135 2.050 4.705 2.210 ;
        RECT 1.135 1.150 1.295 2.050 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 0.175 0.330 2.255 0.490 ;
  END
END OA21D1_2

#--------EOF---------

MACRO OA21D1_3
  CLASS CORE ;
  FOREIGN OA21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 1.390 2.735 2.050 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.945 3.420 4.245 3.720 ;
        RECT 4.030 2.280 4.160 3.420 ;
        RECT 3.945 1.980 4.245 2.280 ;
      LAYER Metal1 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 3.650 4.175 4.630 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 3.965 2.050 4.225 2.210 ;
        RECT 4.015 1.150 4.175 2.050 ;
        RECT 3.965 0.990 4.225 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 4.510 2.760 4.640 4.100 ;
        RECT 4.425 2.460 4.725 2.760 ;
        RECT 4.510 1.620 4.640 2.460 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 4.330 0.335 4.630 ;
        RECT 3.055 4.330 3.215 4.630 ;
        RECT 0.175 4.170 3.215 4.330 ;
        RECT 2.095 2.690 2.255 4.170 ;
        RECT 2.095 2.530 4.705 2.690 ;
        RECT 2.095 1.150 2.255 2.530 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OA21D1_3

#--------EOF---------

MACRO OAI21D1
  CLASS CORE ;
  FOREIGN OAI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.494000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.330 1.295 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 1.150 2.255 4.170 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.150 0.335 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 3.055 4.790 3.215 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OAI21D1

#--------EOF---------

MACRO OAI21D1_1
  CLASS CORE ;
  FOREIGN OAI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.494000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 1.150 1.295 4.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.150 3.215 0.990 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
        RECT 0.175 4.790 0.335 5.970 ;
        RECT 3.055 4.790 3.215 5.970 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 0.175 0.330 2.255 0.490 ;
  END
END OAI21D1_1

#--------EOF---------

MACRO OAI21D1_2
  CLASS CORE ;
  FOREIGN OAI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.034000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.505 4.560 2.805 4.860 ;
        RECT 2.590 1.220 2.720 4.560 ;
        RECT 2.505 0.920 2.805 1.220 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 3.265 4.790 ;
        RECT 0.175 1.150 0.335 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.785 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OAI21D1_2

#--------EOF---------

MACRO OAI21D1_3
  CLASS CORE ;
  FOREIGN OAI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.034000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 4.630 3.265 4.790 ;
        RECT 2.095 1.550 2.255 4.630 ;
        RECT 0.175 1.390 2.255 1.550 ;
        RECT 0.175 1.150 0.335 1.390 ;
        RECT 2.095 1.150 2.255 1.390 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.620 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 2.280 3.680 4.100 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.535 2.210 3.695 2.690 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 1.135 0.330 3.215 0.490 ;
  END
END OAI21D1_3

#--------EOF---------

MACRO OR2D1
  CLASS CORE ;
  FOREIGN OR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.740 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.980275 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 3.240 2.720 4.100 ;
        RECT 2.505 2.940 2.805 3.240 ;
        RECT 2.590 1.555 2.720 2.940 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 3.170 0.335 4.630 ;
        RECT 0.175 3.010 2.785 3.170 ;
        RECT 1.135 1.150 1.295 3.010 ;
        RECT 1.085 0.990 1.345 1.150 ;
  END
END OR2D1

#--------EOF---------

MACRO OR2D1_1
  CLASS CORE ;
  FOREIGN OR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.980275 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 2.505 4.560 2.805 4.860 ;
        RECT 2.590 3.635 2.720 4.560 ;
        RECT 3.550 3.635 3.680 4.100 ;
        RECT 2.590 3.505 3.680 3.635 ;
        RECT 3.550 1.555 3.680 3.505 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 2.785 4.790 ;
        RECT 2.095 4.330 2.255 4.630 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 1.150 1.295 4.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
  END
END OR2D1_1

#--------EOF---------

MACRO OR2D1_2
  CLASS CORE ;
  FOREIGN OR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.980275 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 1.555 3.680 4.100 ;
        RECT 2.025 0.475 2.325 0.560 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 2.025 0.345 3.680 0.475 ;
        RECT 2.025 0.260 2.325 0.345 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 2.255 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 0.125 0.990 2.305 1.150 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 2.045 0.330 2.305 0.490 ;
  END
END OR2D1_2

#--------EOF---------

MACRO OR2D1_3
  CLASS CORE ;
  FOREIGN OR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.420 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.980275 ;
    PORT
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 1.150 3.215 4.630 ;
        RECT 3.005 0.990 3.265 1.150 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 1.630 2.280 1.760 4.100 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.555 1.760 1.980 ;
        RECT 1.630 0.740 1.760 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.210 1.775 2.690 ;
        RECT 1.565 2.050 1.825 2.210 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225550 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.555 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 1.555 3.680 4.100 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 3.465 0.260 3.765 0.560 ;
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 1.150 2.255 4.630 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.175 0.490 0.335 0.990 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 0.175 0.330 3.745 0.490 ;
  END
END OR2D1_3

#--------EOF---------

MACRO TAPCELL
  CLASS CORE ;
  FOREIGN TAPCELL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.380 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.340 0.920 0.600 1.080 ;
        RECT 0.820 0.920 1.080 1.080 ;
        RECT 1.300 0.920 1.560 1.080 ;
        RECT 0.390 0.150 0.550 0.920 ;
        RECT 0.870 0.150 1.030 0.920 ;
        RECT 1.350 0.150 1.510 0.920 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 2.380 6.270 ;
        RECT 0.390 4.860 0.550 5.970 ;
        RECT 0.870 4.860 1.030 5.970 ;
        RECT 1.350 4.860 1.510 5.970 ;
        RECT 0.340 4.700 0.600 4.860 ;
        RECT 0.820 4.700 1.080 4.860 ;
        RECT 1.300 4.700 1.560 4.860 ;
    END
  END vdd
END TAPCELL

#--------EOF---------

MACRO TIEH
  CLASS CORE ;
  FOREIGN TIEH ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 4.790 0.815 5.130 ;
        RECT 0.175 4.630 0.815 4.790 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 1.620 0.800 4.100 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH

#--------EOF---------

MACRO TIEH_1
  CLASS CORE ;
  FOREIGN TIEH_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 4.790 0.815 5.130 ;
        RECT 0.175 4.630 0.815 4.790 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 1.620 0.800 4.100 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH_1

#--------EOF---------

MACRO TIEH_2
  CLASS CORE ;
  FOREIGN TIEH_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 4.790 0.815 5.130 ;
        RECT 0.175 4.630 0.815 4.790 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 1.620 0.800 4.100 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH_2

#--------EOF---------

MACRO TIEH_3
  CLASS CORE ;
  FOREIGN TIEH_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 4.790 0.815 5.130 ;
        RECT 0.175 4.630 0.815 4.790 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 1.620 0.800 4.100 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 0.990 0.815 1.150 ;
        RECT 0.655 0.490 0.815 0.990 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH_3

#--------EOF---------

MACRO TIEL
  CLASS CORE ;
  FOREIGN TIEL ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 1.150 0.815 1.550 ;
        RECT 0.175 0.990 0.815 1.150 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.670 1.620 0.800 3.420 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 0.605 3.490 0.865 3.650 ;
  END
END TIEL

#--------EOF---------

MACRO TIEL_1
  CLASS CORE ;
  FOREIGN TIEL_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 1.150 0.815 1.550 ;
        RECT 0.175 0.990 0.815 1.150 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.670 1.620 0.800 3.420 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 0.605 3.490 0.865 3.650 ;
  END
END TIEL_1

#--------EOF---------

MACRO TIEL_2
  CLASS CORE ;
  FOREIGN TIEL_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 1.150 0.815 1.550 ;
        RECT 0.175 0.990 0.815 1.150 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.670 1.620 0.800 3.420 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 0.605 3.490 0.865 3.650 ;
  END
END TIEL_2

#--------EOF---------

MACRO TIEL_3
  CLASS CORE ;
  FOREIGN TIEL_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.700 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 1.150 0.815 1.550 ;
        RECT 0.175 0.990 0.815 1.150 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.150 1.295 0.990 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 1.700 6.270 ;
        RECT 1.135 4.790 1.295 5.970 ;
        RECT 1.085 4.630 1.345 4.790 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 3.720 0.800 4.100 ;
        RECT 0.585 3.420 0.885 3.720 ;
        RECT 0.670 1.620 0.800 3.420 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.125 4.630 0.815 4.790 ;
        RECT 0.655 3.650 0.815 4.630 ;
        RECT 0.605 3.490 0.865 3.650 ;
  END
END TIEL_3

#--------EOF---------

MACRO XNR2D1
  CLASS CORE ;
  FOREIGN XNR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 4.315 2.720 4.650 ;
        RECT 2.110 4.185 2.720 4.315 ;
        RECT 2.110 2.675 2.240 4.185 ;
        RECT 4.510 3.635 4.640 4.650 ;
        RECT 1.630 2.545 2.240 2.675 ;
        RECT 4.030 3.505 4.640 3.635 ;
        RECT 1.630 1.270 1.760 2.545 ;
        RECT 4.030 2.195 4.160 3.505 ;
        RECT 4.030 2.065 4.640 2.195 ;
        RECT 4.510 1.270 4.640 2.065 ;
        RECT 1.630 0.475 1.760 0.920 ;
        RECT 4.510 0.560 4.640 0.920 ;
        RECT 4.425 0.475 4.725 0.560 ;
        RECT 1.630 0.345 4.725 0.475 ;
        RECT 4.425 0.260 4.725 0.345 ;
      LAYER Metal1 ;
        RECT 4.495 0.490 4.655 1.150 ;
        RECT 4.445 0.330 4.705 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.065 5.775 1.365 5.860 ;
        RECT 1.065 5.645 3.680 5.775 ;
        RECT 1.065 5.560 1.365 5.645 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 6.345 5.560 6.645 5.860 ;
        RECT 6.430 5.200 6.560 5.560 ;
        RECT 1.630 3.240 1.760 4.650 ;
        RECT 2.985 4.100 3.285 4.400 ;
        RECT 1.545 2.940 1.845 3.240 ;
        RECT 2.505 2.940 2.805 3.240 ;
        RECT 2.590 1.270 2.720 2.940 ;
        RECT 3.070 2.280 3.200 4.100 ;
        RECT 2.985 1.980 3.285 2.280 ;
        RECT 3.550 1.270 3.680 4.650 ;
        RECT 4.425 2.675 4.725 2.760 ;
        RECT 6.430 2.675 6.560 4.100 ;
        RECT 4.425 2.545 6.560 2.675 ;
        RECT 4.425 2.460 4.725 2.545 ;
        RECT 6.430 1.620 6.560 2.545 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 2.095 5.630 6.625 5.790 ;
        RECT 1.135 5.130 1.295 5.630 ;
        RECT 2.095 5.130 2.255 5.630 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 3.055 4.330 3.215 4.970 ;
        RECT 3.005 4.170 3.265 4.330 ;
        RECT 4.975 3.170 5.135 4.970 ;
        RECT 1.565 3.010 5.135 3.170 ;
        RECT 2.095 2.530 4.705 2.690 ;
        RECT 2.095 1.150 2.255 2.530 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.055 1.150 3.215 2.050 ;
        RECT 4.975 1.150 5.135 3.010 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
  END
END XNR2D1

#--------EOF---------

MACRO XNR2D1_1
  CLASS CORE ;
  FOREIGN XNR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 3.720 3.680 4.100 ;
        RECT 3.465 3.420 3.765 3.720 ;
        RECT 3.465 1.980 3.765 2.280 ;
        RECT 3.550 1.620 3.680 1.980 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 3.535 2.210 3.695 3.490 ;
        RECT 3.485 2.050 3.745 2.210 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.645 4.640 5.775 ;
        RECT 1.630 5.200 1.760 5.645 ;
        RECT 4.510 5.200 4.640 5.645 ;
        RECT 1.630 4.470 1.760 4.650 ;
        RECT 4.510 4.400 4.640 4.650 ;
        RECT 4.425 4.100 4.725 4.400 ;
        RECT 4.425 2.460 4.725 2.760 ;
        RECT 2.590 1.270 2.720 1.450 ;
        RECT 4.510 1.270 4.640 2.460 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 4.510 0.475 4.640 0.920 ;
        RECT 2.590 0.345 4.640 0.475 ;
      LAYER Metal1 ;
        RECT 4.445 4.170 4.705 4.330 ;
        RECT 4.495 2.690 4.655 4.170 ;
        RECT 4.445 2.530 4.705 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.150 4.175 0.990 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 4.015 5.130 4.175 5.970 ;
        RECT 3.965 4.970 4.225 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.585 5.560 0.885 5.860 ;
        RECT 0.670 5.200 0.800 5.560 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 1.270 0.800 4.650 ;
        RECT 2.590 2.280 2.720 4.650 ;
        RECT 2.985 3.155 3.285 3.240 ;
        RECT 6.430 3.155 6.560 4.100 ;
        RECT 2.985 3.025 6.560 3.155 ;
        RECT 2.985 2.940 3.285 3.025 ;
        RECT 2.505 2.195 2.805 2.280 ;
        RECT 1.630 2.065 2.805 2.195 ;
        RECT 1.630 1.270 1.760 2.065 ;
        RECT 2.505 1.980 2.805 2.065 ;
        RECT 6.430 1.620 6.560 3.025 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 5.630 3.215 5.790 ;
        RECT 3.055 5.130 3.215 5.630 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 2.095 4.790 2.255 4.970 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 3.055 3.170 3.215 4.630 ;
        RECT 3.005 3.010 3.265 3.170 ;
        RECT 3.055 2.690 3.215 3.010 ;
        RECT 2.095 2.530 3.215 2.690 ;
        RECT 2.095 1.150 2.255 2.530 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 1.550 2.735 2.050 ;
        RECT 4.975 1.550 5.135 4.970 ;
        RECT 2.575 1.390 5.135 1.550 ;
        RECT 4.975 1.150 5.135 1.390 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 3.055 0.490 3.215 0.990 ;
        RECT 0.605 0.330 3.215 0.490 ;
  END
END XNR2D1_1

#--------EOF---------

MACRO XNR2D1_2
  CLASS CORE ;
  FOREIGN XNR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 2.050 3.215 2.210 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 1.150 7.055 4.630 ;
        RECT 6.845 0.990 7.105 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 3.155 0.800 4.650 ;
        RECT 1.545 3.155 1.845 3.240 ;
        RECT 0.670 3.025 1.845 3.155 ;
        RECT 1.545 2.940 1.845 3.025 ;
        RECT 2.985 3.155 3.285 3.240 ;
        RECT 3.550 3.155 3.680 4.650 ;
        RECT 2.985 3.025 3.680 3.155 ;
        RECT 2.985 2.940 3.285 3.025 ;
        RECT 1.630 1.270 1.760 2.940 ;
        RECT 3.070 2.195 3.200 2.940 ;
        RECT 3.070 2.065 3.680 2.195 ;
        RECT 3.550 1.270 3.680 2.065 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 1.565 3.010 3.265 3.170 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
        RECT 5.935 5.130 6.095 5.970 ;
        RECT 5.885 4.970 6.145 5.130 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 1.630 3.635 1.760 4.650 ;
        RECT 5.470 4.400 5.600 4.650 ;
        RECT 3.945 4.315 4.245 4.400 ;
        RECT 5.385 4.315 5.685 4.400 ;
        RECT 3.945 4.185 5.685 4.315 ;
        RECT 3.945 4.100 4.245 4.185 ;
        RECT 5.385 4.100 5.685 4.185 ;
        RECT 1.630 3.505 2.240 3.635 ;
        RECT 2.110 2.280 2.240 3.505 ;
        RECT 3.465 2.675 3.765 2.760 ;
        RECT 6.430 2.675 6.560 4.100 ;
        RECT 3.465 2.545 6.560 2.675 ;
        RECT 3.465 2.460 3.765 2.545 ;
        RECT 2.025 1.980 2.325 2.280 ;
        RECT 6.430 1.620 6.560 2.545 ;
        RECT 0.670 1.270 0.800 1.450 ;
        RECT 5.470 1.270 5.600 1.450 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 5.470 0.560 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
        RECT 5.385 0.260 5.685 0.560 ;
      LAYER Metal1 ;
        RECT 0.175 5.630 5.135 5.790 ;
        RECT 0.175 5.130 0.335 5.630 ;
        RECT 4.975 5.130 5.135 5.630 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.965 4.970 4.655 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 1.135 2.690 1.295 4.970 ;
        RECT 2.045 4.630 4.175 4.790 ;
        RECT 4.015 4.330 4.175 4.630 ;
        RECT 3.965 4.170 4.225 4.330 ;
        RECT 1.135 2.530 3.745 2.690 ;
        RECT 1.135 1.150 1.295 2.530 ;
        RECT 2.045 2.050 2.305 2.210 ;
        RECT 2.095 1.550 2.255 2.050 ;
        RECT 4.495 1.550 4.655 4.970 ;
        RECT 1.615 1.390 4.655 1.550 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.615 0.490 1.775 1.390 ;
        RECT 4.015 1.150 4.175 1.390 ;
        RECT 4.975 1.150 5.135 4.970 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.605 0.330 1.775 0.490 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 5.455 0.490 5.615 4.170 ;
        RECT 2.095 0.330 5.665 0.490 ;
  END
END XNR2D1_2

#--------EOF---------

MACRO XNR2D1_3
  CLASS CORE ;
  FOREIGN XNR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 1.150 5.135 4.630 ;
        RECT 4.925 0.990 5.185 1.150 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 0.670 4.400 0.800 4.650 ;
        RECT 3.550 4.400 3.680 4.650 ;
        RECT 0.585 4.100 0.885 4.400 ;
        RECT 3.465 4.100 3.765 4.400 ;
        RECT 1.630 1.270 1.760 1.450 ;
        RECT 3.550 1.270 3.680 4.100 ;
        RECT 1.630 0.560 1.760 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 1.545 0.260 1.845 0.560 ;
        RECT 3.465 0.260 3.765 0.560 ;
      LAYER Metal1 ;
        RECT 0.605 4.170 3.745 4.330 ;
        RECT 1.565 0.330 3.745 0.490 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 4.425 4.900 4.725 5.200 ;
        RECT 1.630 4.470 1.760 4.650 ;
        RECT 4.510 3.635 4.640 4.900 ;
        RECT 5.470 3.920 5.600 4.100 ;
        RECT 5.385 3.635 5.685 3.720 ;
        RECT 4.510 3.505 5.685 3.635 ;
        RECT 5.385 3.420 5.685 3.505 ;
        RECT 5.470 1.620 5.600 1.800 ;
        RECT 0.670 1.270 0.800 1.450 ;
        RECT 6.430 1.270 6.560 4.650 ;
        RECT 0.670 0.740 0.800 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.560 6.560 0.920 ;
        RECT 6.345 0.260 6.645 0.560 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 7.105 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 2.045 4.630 4.175 4.790 ;
        RECT 4.015 1.150 4.175 4.630 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 5.455 1.150 5.615 3.490 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 4.655 1.150 ;
        RECT 5.455 0.990 7.105 1.150 ;
        RECT 4.495 0.490 4.655 0.990 ;
        RECT 4.495 0.330 6.625 0.490 ;
  END
END XNR2D1_3

#--------EOF---------

MACRO XOR2D1
  CLASS CORE ;
  FOREIGN XOR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 2.590 4.400 2.720 4.650 ;
        RECT 4.510 4.400 4.640 4.650 ;
        RECT 2.505 4.100 2.805 4.400 ;
        RECT 4.425 4.100 4.725 4.400 ;
        RECT 4.510 2.760 4.640 4.100 ;
        RECT 1.545 2.460 1.845 2.760 ;
        RECT 4.425 2.460 4.725 2.760 ;
        RECT 1.630 1.270 1.760 2.460 ;
        RECT 4.510 1.270 4.640 2.460 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 4.170 4.705 4.330 ;
        RECT 1.565 2.530 4.705 2.690 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 3.550 3.720 3.680 4.100 ;
        RECT 3.465 3.420 3.765 3.720 ;
        RECT 3.550 1.620 3.680 3.420 ;
        RECT 3.550 0.740 3.680 0.920 ;
      LAYER Metal1 ;
        RECT 3.485 3.490 4.175 3.650 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.585 5.560 0.885 5.860 ;
        RECT 0.670 5.200 0.800 5.560 ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 1.270 0.800 4.650 ;
        RECT 1.630 3.240 1.760 4.650 ;
        RECT 2.025 3.420 2.325 3.720 ;
        RECT 1.545 2.940 1.845 3.240 ;
        RECT 2.110 2.280 2.240 3.420 ;
        RECT 2.505 2.940 2.805 3.240 ;
        RECT 2.025 1.980 2.325 2.280 ;
        RECT 2.590 1.270 2.720 2.940 ;
        RECT 4.905 2.195 5.205 2.280 ;
        RECT 6.430 2.195 6.560 4.100 ;
        RECT 4.905 2.065 6.560 2.195 ;
        RECT 4.905 1.980 5.205 2.065 ;
        RECT 6.430 1.620 6.560 2.065 ;
        RECT 0.670 0.560 0.800 0.920 ;
        RECT 0.585 0.260 0.885 0.560 ;
        RECT 2.590 0.475 2.720 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 2.985 0.475 3.285 0.560 ;
        RECT 2.590 0.345 3.285 0.475 ;
        RECT 2.985 0.260 3.285 0.345 ;
      LAYER Metal1 ;
        RECT 0.605 5.630 3.215 5.790 ;
        RECT 3.055 5.130 3.215 5.630 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.135 1.150 1.295 4.970 ;
        RECT 2.095 3.650 2.255 4.970 ;
        RECT 2.045 3.490 2.305 3.650 ;
        RECT 4.975 3.170 5.135 4.970 ;
        RECT 1.565 3.010 5.135 3.170 ;
        RECT 2.045 2.050 5.185 2.210 ;
        RECT 2.095 1.150 2.255 2.050 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.575 0.990 3.265 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 2.575 0.490 2.735 0.990 ;
        RECT 4.975 0.490 5.135 0.990 ;
        RECT 0.605 0.330 2.735 0.490 ;
        RECT 3.005 0.330 5.135 0.490 ;
  END
END XOR2D1

#--------EOF---------

MACRO XOR2D1_1
  CLASS CORE ;
  FOREIGN XOR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 1.630 4.315 1.760 4.650 ;
        RECT 1.150 4.185 1.760 4.315 ;
        RECT 1.150 3.635 1.280 4.185 ;
        RECT 0.670 3.505 1.280 3.635 ;
        RECT 0.670 1.270 0.800 3.505 ;
        RECT 3.550 1.270 3.680 4.650 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 2.505 0.475 2.805 0.560 ;
        RECT 0.670 0.345 2.805 0.475 ;
        RECT 2.505 0.260 2.805 0.345 ;
        RECT 3.465 0.260 3.765 0.560 ;
      LAYER Metal1 ;
        RECT 2.525 0.330 3.745 0.490 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.525 2.050 3.215 2.210 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 1.150 7.055 4.630 ;
        RECT 6.845 0.990 7.105 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.585 5.560 0.885 5.860 ;
        RECT 0.670 5.200 0.800 5.560 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 4.470 0.800 4.650 ;
        RECT 5.470 4.470 5.600 4.650 ;
        RECT 1.545 3.420 1.845 3.720 ;
        RECT 1.630 2.675 1.760 3.420 ;
        RECT 2.025 2.675 2.325 2.760 ;
        RECT 1.630 2.545 2.325 2.675 ;
        RECT 1.630 1.270 1.760 2.545 ;
        RECT 2.025 2.460 2.325 2.545 ;
        RECT 4.425 2.675 4.725 2.760 ;
        RECT 5.385 2.675 5.685 2.760 ;
        RECT 4.425 2.545 5.685 2.675 ;
        RECT 4.425 2.460 4.725 2.545 ;
        RECT 5.385 2.460 5.685 2.545 ;
        RECT 6.430 2.195 6.560 4.100 ;
        RECT 4.990 2.065 6.560 2.195 ;
        RECT 4.425 1.535 4.725 1.620 ;
        RECT 4.990 1.535 5.120 2.065 ;
        RECT 6.430 1.620 6.560 2.065 ;
        RECT 4.425 1.405 5.120 1.535 ;
        RECT 4.425 1.320 4.725 1.405 ;
        RECT 5.470 1.270 5.600 1.450 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 5.470 0.740 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
      LAYER Metal1 ;
        RECT 0.605 5.630 1.775 5.790 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 1.135 1.550 1.295 4.970 ;
        RECT 1.615 3.650 1.775 5.630 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 4.015 2.690 4.175 4.970 ;
        RECT 2.045 2.530 4.705 2.690 ;
        RECT 1.135 1.390 4.705 1.550 ;
        RECT 1.135 1.150 1.295 1.390 ;
        RECT 4.975 1.150 5.135 4.970 ;
        RECT 5.405 2.530 5.665 2.690 ;
        RECT 0.125 0.990 5.185 1.150 ;
        RECT 4.015 0.490 4.175 0.990 ;
        RECT 5.455 0.490 5.615 2.530 ;
        RECT 4.015 0.330 5.615 0.490 ;
  END
END XOR2D1_1

#--------EOF---------

MACRO XOR2D1_2
  CLASS CORE ;
  FOREIGN XOR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 3.550 5.200 3.680 5.380 ;
        RECT 1.630 4.315 1.760 4.650 ;
        RECT 1.150 4.185 1.760 4.315 ;
        RECT 1.150 3.635 1.280 4.185 ;
        RECT 0.670 3.505 1.280 3.635 ;
        RECT 0.670 1.270 0.800 3.505 ;
        RECT 3.550 1.270 3.680 4.650 ;
        RECT 0.670 0.475 0.800 0.920 ;
        RECT 3.550 0.560 3.680 0.920 ;
        RECT 2.505 0.475 2.805 0.560 ;
        RECT 0.670 0.345 2.805 0.475 ;
        RECT 2.505 0.260 2.805 0.345 ;
        RECT 3.465 0.260 3.765 0.560 ;
      LAYER Metal1 ;
        RECT 2.525 0.330 3.745 0.490 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 2.590 2.280 2.720 4.100 ;
        RECT 2.505 1.980 2.805 2.280 ;
        RECT 2.590 1.620 2.720 1.980 ;
        RECT 2.590 0.740 2.720 0.920 ;
      LAYER Metal1 ;
        RECT 2.575 2.210 2.735 2.690 ;
        RECT 2.525 2.050 2.785 2.210 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 1.150 5.135 4.630 ;
        RECT 4.925 0.990 5.185 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 5.470 5.200 5.600 5.380 ;
        RECT 6.430 5.200 6.560 5.380 ;
        RECT 0.670 4.470 0.800 4.650 ;
        RECT 6.430 4.470 6.560 4.650 ;
        RECT 5.470 1.620 5.600 4.100 ;
        RECT 1.630 1.270 1.760 1.450 ;
        RECT 4.425 1.320 4.725 1.620 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 4.510 0.475 4.640 1.320 ;
        RECT 6.430 1.270 6.560 1.450 ;
        RECT 5.470 0.475 5.600 0.920 ;
        RECT 6.430 0.740 6.560 0.920 ;
        RECT 4.510 0.345 5.600 0.475 ;
      LAYER Metal1 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 0.175 1.150 0.335 4.970 ;
        RECT 1.135 1.550 1.295 4.970 ;
        RECT 1.135 1.390 4.705 1.550 ;
        RECT 1.135 1.150 1.295 1.390 ;
        RECT 6.895 1.150 7.055 4.970 ;
        RECT 0.125 0.990 4.655 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 4.495 0.490 4.655 0.990 ;
        RECT 6.895 0.490 7.055 0.990 ;
        RECT 4.495 0.330 7.055 0.490 ;
  END
END XOR2D1_2

#--------EOF---------

MACRO XOR2D1_3
  CLASS CORE ;
  FOREIGN XOR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.630 5.200 1.760 5.380 ;
        RECT 4.510 5.200 4.640 5.380 ;
        RECT 1.630 2.760 1.760 4.650 ;
        RECT 1.545 2.675 1.845 2.760 ;
        RECT 1.545 2.545 2.720 2.675 ;
        RECT 1.545 2.460 1.845 2.545 ;
        RECT 2.590 2.195 2.720 2.545 ;
        RECT 4.510 2.195 4.640 4.650 ;
        RECT 2.590 2.065 4.640 2.195 ;
        RECT 2.590 1.270 2.720 2.065 ;
        RECT 4.510 1.270 4.640 2.065 ;
        RECT 2.590 0.740 2.720 0.920 ;
        RECT 4.510 0.740 4.640 0.920 ;
      LAYER Metal1 ;
        RECT 1.615 2.690 1.775 3.170 ;
        RECT 1.565 2.530 1.825 2.690 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.234000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.670 5.200 0.800 5.380 ;
        RECT 0.670 2.280 0.800 4.100 ;
        RECT 0.585 1.980 0.885 2.280 ;
        RECT 0.670 1.620 0.800 1.980 ;
        RECT 0.670 0.740 0.800 0.920 ;
      LAYER Metal1 ;
        RECT 0.655 2.210 0.815 2.690 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.017000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 1.150 6.095 4.630 ;
        RECT 5.885 0.990 6.145 1.150 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END
  END vdd
  OBS
      LAYER GatPoly ;
        RECT 1.065 5.775 1.365 5.860 ;
        RECT 1.065 5.645 3.680 5.775 ;
        RECT 1.065 5.560 1.365 5.645 ;
        RECT 2.590 5.200 2.720 5.380 ;
        RECT 3.550 5.200 3.680 5.645 ;
        RECT 6.345 5.560 6.645 5.860 ;
        RECT 6.430 5.200 6.560 5.560 ;
        RECT 2.590 3.240 2.720 4.650 ;
        RECT 3.550 4.470 3.680 4.650 ;
        RECT 2.505 3.155 2.805 3.240 ;
        RECT 3.945 3.155 4.245 3.240 ;
        RECT 2.505 3.025 4.245 3.155 ;
        RECT 2.505 2.940 2.805 3.025 ;
        RECT 3.945 2.940 4.245 3.025 ;
        RECT 1.545 1.980 1.845 2.280 ;
        RECT 1.630 1.270 1.760 1.980 ;
        RECT 6.430 1.620 6.560 4.100 ;
        RECT 3.550 1.270 3.680 1.450 ;
        RECT 1.630 0.740 1.760 0.920 ;
        RECT 1.065 0.475 1.365 0.560 ;
        RECT 3.550 0.475 3.680 0.920 ;
        RECT 6.430 0.560 6.560 0.920 ;
        RECT 1.065 0.345 3.680 0.475 ;
        RECT 1.065 0.260 1.365 0.345 ;
        RECT 6.345 0.260 6.645 0.560 ;
      LAYER Metal1 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 2.095 5.630 6.625 5.790 ;
        RECT 1.135 5.130 1.295 5.630 ;
        RECT 2.095 5.130 2.255 5.630 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 4.970 3.695 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 1.150 1.295 4.630 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 2.575 2.210 2.735 3.010 ;
        RECT 1.565 2.050 2.735 2.210 ;
        RECT 3.535 1.150 3.695 4.970 ;
        RECT 4.975 4.790 5.135 4.970 ;
        RECT 4.015 4.630 5.135 4.790 ;
        RECT 4.015 3.170 4.175 4.630 ;
        RECT 3.965 3.010 4.225 3.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.695 1.150 ;
        RECT 4.015 1.150 4.175 3.010 ;
        RECT 4.015 0.990 5.185 1.150 ;
        RECT 1.135 0.490 1.295 0.990 ;
        RECT 2.095 0.490 2.255 0.990 ;
        RECT 1.085 0.330 1.345 0.490 ;
        RECT 2.095 0.330 6.625 0.490 ;
  END
END XOR2D1_3

#--------EOF---------


END LIBRARY
