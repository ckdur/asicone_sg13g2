VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MACRO sg13g2_bpd60
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd60 0 0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 67.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 62.930 60.000 67.000 ;
        RECT 0.000 11.070 4.070 62.930 ;
        RECT 55.930 11.070 60.000 62.930 ;
        RECT 0.000 7.000 60.000 11.070 ;
        RECT 6.500 0.000 13.500 7.000 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
      LAYER Metal4 ;
        RECT 0.000 62.930 60.000 67.000 ;
        RECT 0.000 11.070 4.070 62.930 ;
        RECT 55.930 11.070 60.000 62.930 ;
        RECT 0.000 7.000 60.000 11.070 ;
        RECT 6.500 0.000 13.500 7.000 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
      LAYER Metal5 ;
        RECT 0.000 62.930 60.000 67.000 ;
        RECT 0.000 11.070 4.070 62.930 ;
        RECT 55.930 11.070 60.000 62.930 ;
        RECT 0.000 7.000 60.000 11.070 ;
        RECT 6.500 0.000 13.500 7.000 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
      LAYER TopMetal1 ;
        RECT 0.000 62.930 60.000 67.000 ;
        RECT 0.000 11.070 4.070 62.930 ;
        RECT 55.930 11.070 60.000 62.930 ;
        RECT 0.000 7.000 60.000 11.070 ;
        RECT 6.500 0.000 13.500 7.000 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 64.900 60.000 67.000 ;
        RECT 0.000 64.015 2.985 64.900 ;
        RECT 3.080 64.015 4.980 64.900 ;
        RECT 5.080 64.015 6.980 64.900 ;
        RECT 7.075 64.015 8.975 64.900 ;
        RECT 9.075 64.015 10.975 64.900 ;
        RECT 11.070 64.015 12.970 64.900 ;
        RECT 13.070 64.015 14.970 64.900 ;
        RECT 15.065 64.015 16.965 64.900 ;
        RECT 17.065 64.015 18.965 64.900 ;
        RECT 19.060 64.015 20.960 64.900 ;
        RECT 21.060 64.015 22.960 64.900 ;
        RECT 23.055 64.015 24.955 64.900 ;
        RECT 25.055 64.015 26.955 64.900 ;
        RECT 27.050 64.015 28.950 64.900 ;
        RECT 29.050 64.015 30.950 64.900 ;
        RECT 31.045 64.015 32.945 64.900 ;
        RECT 33.045 64.015 34.945 64.900 ;
        RECT 35.040 64.015 36.940 64.900 ;
        RECT 37.040 64.015 38.940 64.900 ;
        RECT 39.035 64.015 40.935 64.900 ;
        RECT 41.035 64.015 42.935 64.900 ;
        RECT 43.030 64.015 44.930 64.900 ;
        RECT 45.030 64.015 46.930 64.900 ;
        RECT 47.025 64.015 48.925 64.900 ;
        RECT 49.025 64.015 50.925 64.900 ;
        RECT 51.020 64.015 52.920 64.900 ;
        RECT 53.020 64.015 54.920 64.900 ;
        RECT 55.015 64.015 56.915 64.900 ;
        RECT 57.015 64.015 60.000 64.900 ;
        RECT 0.000 63.945 2.100 64.015 ;
        RECT 57.900 63.945 60.000 64.015 ;
        RECT 0.000 62.045 2.985 63.945 ;
        RECT 57.015 62.045 60.000 63.945 ;
        RECT 0.000 61.945 2.100 62.045 ;
        RECT 57.900 61.945 60.000 62.045 ;
        RECT 0.000 60.045 2.985 61.945 ;
        RECT 57.015 60.045 60.000 61.945 ;
        RECT 0.000 59.945 2.100 60.045 ;
        RECT 57.900 59.945 60.000 60.045 ;
        RECT 0.000 58.045 2.985 59.945 ;
        RECT 57.015 58.045 60.000 59.945 ;
        RECT 0.000 57.945 2.100 58.045 ;
        RECT 57.900 57.945 60.000 58.045 ;
        RECT 0.000 56.045 2.985 57.945 ;
        RECT 57.015 56.045 60.000 57.945 ;
        RECT 0.000 55.945 2.100 56.045 ;
        RECT 57.900 55.945 60.000 56.045 ;
        RECT 0.000 54.045 2.985 55.945 ;
        RECT 57.015 54.045 60.000 55.945 ;
        RECT 0.000 53.945 2.100 54.045 ;
        RECT 57.900 53.945 60.000 54.045 ;
        RECT 0.000 52.045 2.985 53.945 ;
        RECT 57.015 52.045 60.000 53.945 ;
        RECT 0.000 51.945 2.100 52.045 ;
        RECT 57.900 51.945 60.000 52.045 ;
        RECT 0.000 50.045 2.985 51.945 ;
        RECT 57.015 50.045 60.000 51.945 ;
        RECT 0.000 49.945 2.100 50.045 ;
        RECT 57.900 49.945 60.000 50.045 ;
        RECT 0.000 48.045 2.985 49.945 ;
        RECT 57.015 48.045 60.000 49.945 ;
        RECT 0.000 47.945 2.100 48.045 ;
        RECT 57.900 47.945 60.000 48.045 ;
        RECT 0.000 46.045 2.985 47.945 ;
        RECT 57.015 46.045 60.000 47.945 ;
        RECT 0.000 45.945 2.100 46.045 ;
        RECT 57.900 45.945 60.000 46.045 ;
        RECT 0.000 44.045 2.985 45.945 ;
        RECT 57.015 44.045 60.000 45.945 ;
        RECT 0.000 43.945 2.100 44.045 ;
        RECT 57.900 43.945 60.000 44.045 ;
        RECT 0.000 42.045 2.985 43.945 ;
        RECT 57.015 42.045 60.000 43.945 ;
        RECT 0.000 41.945 2.100 42.045 ;
        RECT 57.900 41.945 60.000 42.045 ;
        RECT 0.000 40.045 2.985 41.945 ;
        RECT 57.015 40.045 60.000 41.945 ;
        RECT 0.000 39.945 2.100 40.045 ;
        RECT 57.900 39.945 60.000 40.045 ;
        RECT 0.000 38.045 2.985 39.945 ;
        RECT 57.015 38.045 60.000 39.945 ;
        RECT 0.000 37.950 2.100 38.045 ;
        RECT 57.900 37.950 60.000 38.045 ;
        RECT 0.000 36.050 2.985 37.950 ;
        RECT 57.015 36.050 60.000 37.950 ;
        RECT 0.000 35.950 2.100 36.050 ;
        RECT 57.900 35.950 60.000 36.050 ;
        RECT 0.000 34.050 2.985 35.950 ;
        RECT 57.015 34.050 60.000 35.950 ;
        RECT 0.000 33.950 2.100 34.050 ;
        RECT 57.900 33.950 60.000 34.050 ;
        RECT 0.000 32.050 2.985 33.950 ;
        RECT 57.015 32.050 60.000 33.950 ;
        RECT 0.000 31.950 2.100 32.050 ;
        RECT 57.900 31.950 60.000 32.050 ;
        RECT 0.000 30.050 2.985 31.950 ;
        RECT 57.015 30.050 60.000 31.950 ;
        RECT 0.000 29.950 2.100 30.050 ;
        RECT 57.900 29.950 60.000 30.050 ;
        RECT 0.000 28.050 2.985 29.950 ;
        RECT 57.015 28.050 60.000 29.950 ;
        RECT 0.000 27.950 2.100 28.050 ;
        RECT 57.900 27.950 60.000 28.050 ;
        RECT 0.000 26.050 2.985 27.950 ;
        RECT 57.015 26.050 60.000 27.950 ;
        RECT 0.000 25.950 2.100 26.050 ;
        RECT 57.900 25.950 60.000 26.050 ;
        RECT 0.000 24.050 2.985 25.950 ;
        RECT 57.015 24.050 60.000 25.950 ;
        RECT 0.000 23.950 2.100 24.050 ;
        RECT 57.900 23.950 60.000 24.050 ;
        RECT 0.000 22.050 2.985 23.950 ;
        RECT 57.015 22.050 60.000 23.950 ;
        RECT 0.000 21.950 2.100 22.050 ;
        RECT 57.900 21.950 60.000 22.050 ;
        RECT 0.000 20.050 2.985 21.950 ;
        RECT 57.015 20.050 60.000 21.950 ;
        RECT 0.000 19.950 2.100 20.050 ;
        RECT 57.900 19.950 60.000 20.050 ;
        RECT 0.000 18.050 2.985 19.950 ;
        RECT 57.015 18.050 60.000 19.950 ;
        RECT 0.000 17.950 2.100 18.050 ;
        RECT 57.900 17.950 60.000 18.050 ;
        RECT 0.000 16.050 2.985 17.950 ;
        RECT 57.015 16.050 60.000 17.950 ;
        RECT 0.000 15.950 2.100 16.050 ;
        RECT 57.900 15.950 60.000 16.050 ;
        RECT 0.000 14.050 2.985 15.950 ;
        RECT 57.015 14.050 60.000 15.950 ;
        RECT 0.000 13.950 2.100 14.050 ;
        RECT 57.900 13.950 60.000 14.050 ;
        RECT 0.000 12.050 2.985 13.950 ;
        RECT 57.015 12.050 60.000 13.950 ;
        RECT 0.000 11.955 2.100 12.050 ;
        RECT 57.900 11.955 60.000 12.050 ;
        RECT 0.000 10.055 2.985 11.955 ;
        RECT 57.015 10.055 60.000 11.955 ;
        RECT 0.000 9.985 2.100 10.055 ;
        RECT 57.900 9.985 60.000 10.055 ;
        RECT 0.000 9.100 2.985 9.985 ;
        RECT 3.080 9.100 4.980 9.985 ;
        RECT 5.080 9.100 6.980 9.985 ;
        RECT 7.075 9.100 8.975 9.985 ;
        RECT 9.075 9.100 10.975 9.985 ;
        RECT 11.070 9.100 12.970 9.985 ;
        RECT 13.070 9.100 14.970 9.985 ;
        RECT 15.065 9.100 16.965 9.985 ;
        RECT 17.065 9.100 18.965 9.985 ;
        RECT 19.060 9.100 20.960 9.985 ;
        RECT 21.060 9.100 22.960 9.985 ;
        RECT 23.055 9.100 24.955 9.985 ;
        RECT 25.055 9.100 26.955 9.985 ;
        RECT 27.050 9.100 28.950 9.985 ;
        RECT 29.050 9.100 30.950 9.985 ;
        RECT 31.045 9.100 32.945 9.985 ;
        RECT 33.045 9.100 34.945 9.985 ;
        RECT 35.040 9.100 36.940 9.985 ;
        RECT 37.040 9.100 38.940 9.985 ;
        RECT 39.035 9.100 40.935 9.985 ;
        RECT 41.035 9.100 42.935 9.985 ;
        RECT 43.030 9.100 44.930 9.985 ;
        RECT 45.030 9.100 46.930 9.985 ;
        RECT 47.025 9.100 48.925 9.985 ;
        RECT 49.025 9.100 50.925 9.985 ;
        RECT 51.020 9.100 52.920 9.985 ;
        RECT 53.020 9.100 54.920 9.985 ;
        RECT 55.015 9.100 56.915 9.985 ;
        RECT 57.015 9.100 60.000 9.985 ;
        RECT 0.000 7.000 60.000 9.100 ;
        RECT 6.500 0.000 13.500 7.000 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
  END
END sg13g2_bpd60

#--------EOF---------

MACRO sg13g2_bpd70
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd70 0 0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 77.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 72.930 70.000 77.000 ;
        RECT 0.000 11.070 4.070 72.930 ;
        RECT 65.930 11.070 70.000 72.930 ;
        RECT 0.000 7.000 70.000 11.070 ;
        RECT 11.500 0.000 18.500 7.000 ;
        RECT 21.500 0.000 28.500 7.000 ;
        RECT 31.500 0.000 38.500 7.000 ;
        RECT 41.500 0.000 48.500 7.000 ;
        RECT 51.500 0.000 58.500 7.000 ;
      LAYER Metal4 ;
        RECT 0.000 72.930 70.000 77.000 ;
        RECT 0.000 11.070 4.070 72.930 ;
        RECT 65.930 11.070 70.000 72.930 ;
        RECT 0.000 7.000 70.000 11.070 ;
        RECT 11.500 0.000 18.500 7.000 ;
        RECT 21.500 0.000 28.500 7.000 ;
        RECT 31.500 0.000 38.500 7.000 ;
        RECT 41.500 0.000 48.500 7.000 ;
        RECT 51.500 0.000 58.500 7.000 ;
      LAYER Metal5 ;
        RECT 0.000 72.930 70.000 77.000 ;
        RECT 0.000 11.070 4.070 72.930 ;
        RECT 65.930 11.070 70.000 72.930 ;
        RECT 0.000 7.000 70.000 11.070 ;
        RECT 11.500 0.000 18.500 7.000 ;
        RECT 21.500 0.000 28.500 7.000 ;
        RECT 31.500 0.000 38.500 7.000 ;
        RECT 41.500 0.000 48.500 7.000 ;
        RECT 51.500 0.000 58.500 7.000 ;
      LAYER TopMetal1 ;
        RECT 0.000 72.930 70.000 77.000 ;
        RECT 0.000 11.070 4.070 72.930 ;
        RECT 65.930 11.070 70.000 72.930 ;
        RECT 0.000 7.000 70.000 11.070 ;
        RECT 11.500 0.000 18.500 7.000 ;
        RECT 21.500 0.000 28.500 7.000 ;
        RECT 31.500 0.000 38.500 7.000 ;
        RECT 41.500 0.000 48.500 7.000 ;
        RECT 51.500 0.000 58.500 7.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 74.900 70.000 77.000 ;
        RECT 0.000 74.015 2.985 74.900 ;
        RECT 3.080 74.015 4.980 74.900 ;
        RECT 5.080 74.015 6.980 74.900 ;
        RECT 7.075 74.015 8.975 74.900 ;
        RECT 9.075 74.015 10.975 74.900 ;
        RECT 11.070 74.015 12.970 74.900 ;
        RECT 13.070 74.015 14.970 74.900 ;
        RECT 15.070 74.015 16.970 74.900 ;
        RECT 17.065 74.015 18.965 74.900 ;
        RECT 19.065 74.015 20.965 74.900 ;
        RECT 21.060 74.015 22.960 74.900 ;
        RECT 23.060 74.015 24.960 74.900 ;
        RECT 25.055 74.015 26.955 74.900 ;
        RECT 27.055 74.015 28.955 74.900 ;
        RECT 29.055 74.015 30.955 74.900 ;
        RECT 31.050 74.015 32.950 74.900 ;
        RECT 33.050 74.015 34.950 74.900 ;
        RECT 35.045 74.015 36.945 74.900 ;
        RECT 37.045 74.015 38.945 74.900 ;
        RECT 39.040 74.015 40.940 74.900 ;
        RECT 41.040 74.015 42.940 74.900 ;
        RECT 43.040 74.015 44.940 74.900 ;
        RECT 45.035 74.015 46.935 74.900 ;
        RECT 47.035 74.015 48.935 74.900 ;
        RECT 49.030 74.015 50.930 74.900 ;
        RECT 51.030 74.015 52.930 74.900 ;
        RECT 53.025 74.015 54.925 74.900 ;
        RECT 55.025 74.015 56.925 74.900 ;
        RECT 57.025 74.015 58.925 74.900 ;
        RECT 59.020 74.015 60.920 74.900 ;
        RECT 61.020 74.015 62.920 74.900 ;
        RECT 63.015 74.015 64.915 74.900 ;
        RECT 65.015 74.015 66.915 74.900 ;
        RECT 67.015 74.015 70.000 74.900 ;
        RECT 0.000 73.945 2.100 74.015 ;
        RECT 67.900 73.945 70.000 74.015 ;
        RECT 0.000 72.045 2.985 73.945 ;
        RECT 67.015 72.045 70.000 73.945 ;
        RECT 0.000 71.945 2.100 72.045 ;
        RECT 67.900 71.945 70.000 72.045 ;
        RECT 0.000 70.045 2.985 71.945 ;
        RECT 67.015 70.045 70.000 71.945 ;
        RECT 0.000 69.945 2.100 70.045 ;
        RECT 67.900 69.945 70.000 70.045 ;
        RECT 0.000 68.045 2.985 69.945 ;
        RECT 67.015 68.045 70.000 69.945 ;
        RECT 0.000 67.945 2.100 68.045 ;
        RECT 67.900 67.945 70.000 68.045 ;
        RECT 0.000 66.045 2.985 67.945 ;
        RECT 67.015 66.045 70.000 67.945 ;
        RECT 0.000 65.945 2.100 66.045 ;
        RECT 67.900 65.945 70.000 66.045 ;
        RECT 0.000 64.045 2.985 65.945 ;
        RECT 67.015 64.045 70.000 65.945 ;
        RECT 0.000 63.945 2.100 64.045 ;
        RECT 67.900 63.945 70.000 64.045 ;
        RECT 0.000 62.045 2.985 63.945 ;
        RECT 67.015 62.045 70.000 63.945 ;
        RECT 0.000 61.945 2.100 62.045 ;
        RECT 67.900 61.945 70.000 62.045 ;
        RECT 0.000 60.045 2.985 61.945 ;
        RECT 67.015 60.045 70.000 61.945 ;
        RECT 0.000 59.945 2.100 60.045 ;
        RECT 67.900 59.945 70.000 60.045 ;
        RECT 0.000 58.045 2.985 59.945 ;
        RECT 67.015 58.045 70.000 59.945 ;
        RECT 0.000 57.945 2.100 58.045 ;
        RECT 67.900 57.945 70.000 58.045 ;
        RECT 0.000 56.045 2.985 57.945 ;
        RECT 67.015 56.045 70.000 57.945 ;
        RECT 0.000 55.945 2.100 56.045 ;
        RECT 67.900 55.945 70.000 56.045 ;
        RECT 0.000 54.045 2.985 55.945 ;
        RECT 67.015 54.045 70.000 55.945 ;
        RECT 0.000 53.945 2.100 54.045 ;
        RECT 67.900 53.945 70.000 54.045 ;
        RECT 0.000 52.045 2.985 53.945 ;
        RECT 67.015 52.045 70.000 53.945 ;
        RECT 0.000 51.945 2.100 52.045 ;
        RECT 67.900 51.945 70.000 52.045 ;
        RECT 0.000 50.045 2.985 51.945 ;
        RECT 67.015 50.045 70.000 51.945 ;
        RECT 0.000 49.945 2.100 50.045 ;
        RECT 67.900 49.945 70.000 50.045 ;
        RECT 0.000 48.045 2.985 49.945 ;
        RECT 67.015 48.045 70.000 49.945 ;
        RECT 0.000 47.945 2.100 48.045 ;
        RECT 67.900 47.945 70.000 48.045 ;
        RECT 0.000 46.045 2.985 47.945 ;
        RECT 67.015 46.045 70.000 47.945 ;
        RECT 0.000 45.945 2.100 46.045 ;
        RECT 67.900 45.945 70.000 46.045 ;
        RECT 0.000 44.045 2.985 45.945 ;
        RECT 67.015 44.045 70.000 45.945 ;
        RECT 0.000 43.945 2.100 44.045 ;
        RECT 67.900 43.945 70.000 44.045 ;
        RECT 0.000 42.045 2.985 43.945 ;
        RECT 67.015 42.045 70.000 43.945 ;
        RECT 0.000 41.950 2.100 42.045 ;
        RECT 67.900 41.950 70.000 42.045 ;
        RECT 0.000 40.050 2.985 41.950 ;
        RECT 67.015 40.050 70.000 41.950 ;
        RECT 0.000 39.950 2.100 40.050 ;
        RECT 67.900 39.950 70.000 40.050 ;
        RECT 0.000 38.050 2.985 39.950 ;
        RECT 67.015 38.050 70.000 39.950 ;
        RECT 0.000 37.950 2.100 38.050 ;
        RECT 67.900 37.950 70.000 38.050 ;
        RECT 0.000 36.050 2.985 37.950 ;
        RECT 67.015 36.050 70.000 37.950 ;
        RECT 0.000 35.950 2.100 36.050 ;
        RECT 67.900 35.950 70.000 36.050 ;
        RECT 0.000 34.050 2.985 35.950 ;
        RECT 67.015 34.050 70.000 35.950 ;
        RECT 0.000 33.950 2.100 34.050 ;
        RECT 67.900 33.950 70.000 34.050 ;
        RECT 0.000 32.050 2.985 33.950 ;
        RECT 67.015 32.050 70.000 33.950 ;
        RECT 0.000 31.950 2.100 32.050 ;
        RECT 67.900 31.950 70.000 32.050 ;
        RECT 0.000 30.050 2.985 31.950 ;
        RECT 67.015 30.050 70.000 31.950 ;
        RECT 0.000 29.950 2.100 30.050 ;
        RECT 67.900 29.950 70.000 30.050 ;
        RECT 0.000 28.050 2.985 29.950 ;
        RECT 67.015 28.050 70.000 29.950 ;
        RECT 0.000 27.950 2.100 28.050 ;
        RECT 67.900 27.950 70.000 28.050 ;
        RECT 0.000 26.050 2.985 27.950 ;
        RECT 67.015 26.050 70.000 27.950 ;
        RECT 0.000 25.950 2.100 26.050 ;
        RECT 67.900 25.950 70.000 26.050 ;
        RECT 0.000 24.050 2.985 25.950 ;
        RECT 67.015 24.050 70.000 25.950 ;
        RECT 0.000 23.950 2.100 24.050 ;
        RECT 67.900 23.950 70.000 24.050 ;
        RECT 0.000 22.050 2.985 23.950 ;
        RECT 67.015 22.050 70.000 23.950 ;
        RECT 0.000 21.950 2.100 22.050 ;
        RECT 67.900 21.950 70.000 22.050 ;
        RECT 0.000 20.050 2.985 21.950 ;
        RECT 67.015 20.050 70.000 21.950 ;
        RECT 0.000 19.950 2.100 20.050 ;
        RECT 67.900 19.950 70.000 20.050 ;
        RECT 0.000 18.050 2.985 19.950 ;
        RECT 67.015 18.050 70.000 19.950 ;
        RECT 0.000 17.950 2.100 18.050 ;
        RECT 67.900 17.950 70.000 18.050 ;
        RECT 0.000 16.050 2.985 17.950 ;
        RECT 67.015 16.050 70.000 17.950 ;
        RECT 0.000 15.950 2.100 16.050 ;
        RECT 67.900 15.950 70.000 16.050 ;
        RECT 0.000 14.050 2.985 15.950 ;
        RECT 67.015 14.050 70.000 15.950 ;
        RECT 0.000 13.950 2.100 14.050 ;
        RECT 67.900 13.950 70.000 14.050 ;
        RECT 0.000 12.050 2.985 13.950 ;
        RECT 67.015 12.050 70.000 13.950 ;
        RECT 0.000 11.955 2.100 12.050 ;
        RECT 67.900 11.955 70.000 12.050 ;
        RECT 0.000 10.055 2.985 11.955 ;
        RECT 67.015 10.055 70.000 11.955 ;
        RECT 0.000 9.985 2.100 10.055 ;
        RECT 67.900 9.985 70.000 10.055 ;
        RECT 0.000 9.100 2.985 9.985 ;
        RECT 3.080 9.100 4.980 9.985 ;
        RECT 5.080 9.100 6.980 9.985 ;
        RECT 7.075 9.100 8.975 9.985 ;
        RECT 9.075 9.100 10.975 9.985 ;
        RECT 11.070 9.100 12.970 9.985 ;
        RECT 13.070 9.100 14.970 9.985 ;
        RECT 15.070 9.100 16.970 9.985 ;
        RECT 17.065 9.100 18.965 9.985 ;
        RECT 19.065 9.100 20.965 9.985 ;
        RECT 21.060 9.100 22.960 9.985 ;
        RECT 23.060 9.100 24.960 9.985 ;
        RECT 25.055 9.100 26.955 9.985 ;
        RECT 27.055 9.100 28.955 9.985 ;
        RECT 29.055 9.100 30.955 9.985 ;
        RECT 31.050 9.100 32.950 9.985 ;
        RECT 33.050 9.100 34.950 9.985 ;
        RECT 35.045 9.100 36.945 9.985 ;
        RECT 37.045 9.100 38.945 9.985 ;
        RECT 39.040 9.100 40.940 9.985 ;
        RECT 41.040 9.100 42.940 9.985 ;
        RECT 43.040 9.100 44.940 9.985 ;
        RECT 45.035 9.100 46.935 9.985 ;
        RECT 47.035 9.100 48.935 9.985 ;
        RECT 49.030 9.100 50.930 9.985 ;
        RECT 51.030 9.100 52.930 9.985 ;
        RECT 53.025 9.100 54.925 9.985 ;
        RECT 55.025 9.100 56.925 9.985 ;
        RECT 57.025 9.100 58.925 9.985 ;
        RECT 59.020 9.100 60.920 9.985 ;
        RECT 61.020 9.100 62.920 9.985 ;
        RECT 63.015 9.100 64.915 9.985 ;
        RECT 65.015 9.100 66.915 9.985 ;
        RECT 67.015 9.100 70.000 9.985 ;
        RECT 0.000 7.000 70.000 9.100 ;
        RECT 11.500 0.000 18.500 7.000 ;
        RECT 21.500 0.000 28.500 7.000 ;
        RECT 31.500 0.000 38.500 7.000 ;
        RECT 41.500 0.000 48.500 7.000 ;
        RECT 51.500 0.000 58.500 7.000 ;
  END
END sg13g2_bpd70

#--------EOF---------

MACRO sg13g2_bpd80
  CLASS BLOCK ;
  FOREIGN sg13g2_bpd80 0 0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 87.000 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER Metal3 ;
        RECT 0.000 82.930 80.000 87.000 ;
        RECT 0.000 11.070 4.070 82.930 ;
        RECT 75.930 11.070 80.000 82.930 ;
        RECT 0.000 7.000 80.000 11.070 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
        RECT 56.500 0.000 63.500 7.000 ;
      LAYER Metal4 ;
        RECT 0.000 82.930 80.000 87.000 ;
        RECT 0.000 11.070 4.070 82.930 ;
        RECT 75.930 11.070 80.000 82.930 ;
        RECT 0.000 7.000 80.000 11.070 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
        RECT 56.500 0.000 63.500 7.000 ;
      LAYER Metal5 ;
        RECT 0.000 82.930 80.000 87.000 ;
        RECT 0.000 11.070 4.070 82.930 ;
        RECT 75.930 11.070 80.000 82.930 ;
        RECT 0.000 7.000 80.000 11.070 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
        RECT 56.500 0.000 63.500 7.000 ;
      LAYER TopMetal1 ;
        RECT 0.000 82.930 80.000 87.000 ;
        RECT 0.000 11.070 4.070 82.930 ;
        RECT 75.930 11.070 80.000 82.930 ;
        RECT 0.000 7.000 80.000 11.070 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
        RECT 56.500 0.000 63.500 7.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 84.900 80.000 87.000 ;
        RECT 0.000 84.015 2.985 84.900 ;
        RECT 3.080 84.015 4.980 84.900 ;
        RECT 5.080 84.015 6.980 84.900 ;
        RECT 7.075 84.015 8.975 84.900 ;
        RECT 9.075 84.015 10.975 84.900 ;
        RECT 11.075 84.015 12.975 84.900 ;
        RECT 13.070 84.015 14.970 84.900 ;
        RECT 15.070 84.015 16.970 84.900 ;
        RECT 17.070 84.015 18.970 84.900 ;
        RECT 19.065 84.015 20.965 84.900 ;
        RECT 21.065 84.015 22.965 84.900 ;
        RECT 23.060 84.015 24.960 84.900 ;
        RECT 25.060 84.015 26.960 84.900 ;
        RECT 27.060 84.015 28.960 84.900 ;
        RECT 29.055 84.015 30.955 84.900 ;
        RECT 31.055 84.015 32.955 84.900 ;
        RECT 33.055 84.015 34.955 84.900 ;
        RECT 35.050 84.015 36.950 84.900 ;
        RECT 37.050 84.015 38.950 84.900 ;
        RECT 39.050 84.015 40.950 84.900 ;
        RECT 41.045 84.015 42.945 84.900 ;
        RECT 43.045 84.015 44.945 84.900 ;
        RECT 45.040 84.015 46.940 84.900 ;
        RECT 47.040 84.015 48.940 84.900 ;
        RECT 49.040 84.015 50.940 84.900 ;
        RECT 51.035 84.015 52.935 84.900 ;
        RECT 53.035 84.015 54.935 84.900 ;
        RECT 55.035 84.015 56.935 84.900 ;
        RECT 57.030 84.015 58.930 84.900 ;
        RECT 59.030 84.015 60.930 84.900 ;
        RECT 61.025 84.015 62.925 84.900 ;
        RECT 63.025 84.015 64.925 84.900 ;
        RECT 65.025 84.015 66.925 84.900 ;
        RECT 67.020 84.015 68.920 84.900 ;
        RECT 69.020 84.015 70.920 84.900 ;
        RECT 71.020 84.015 72.920 84.900 ;
        RECT 73.015 84.015 74.915 84.900 ;
        RECT 75.015 84.015 76.915 84.900 ;
        RECT 77.015 84.015 80.000 84.900 ;
        RECT 0.000 83.945 2.100 84.015 ;
        RECT 77.900 83.945 80.000 84.015 ;
        RECT 0.000 82.045 2.985 83.945 ;
        RECT 77.015 82.045 80.000 83.945 ;
        RECT 0.000 81.945 2.100 82.045 ;
        RECT 77.900 81.945 80.000 82.045 ;
        RECT 0.000 80.045 2.985 81.945 ;
        RECT 77.015 80.045 80.000 81.945 ;
        RECT 0.000 79.945 2.100 80.045 ;
        RECT 77.900 79.945 80.000 80.045 ;
        RECT 0.000 78.045 2.985 79.945 ;
        RECT 77.015 78.045 80.000 79.945 ;
        RECT 0.000 77.945 2.100 78.045 ;
        RECT 77.900 77.945 80.000 78.045 ;
        RECT 0.000 76.045 2.985 77.945 ;
        RECT 77.015 76.045 80.000 77.945 ;
        RECT 0.000 75.945 2.100 76.045 ;
        RECT 77.900 75.945 80.000 76.045 ;
        RECT 0.000 74.045 2.985 75.945 ;
        RECT 77.015 74.045 80.000 75.945 ;
        RECT 0.000 73.945 2.100 74.045 ;
        RECT 77.900 73.945 80.000 74.045 ;
        RECT 0.000 72.045 2.985 73.945 ;
        RECT 77.015 72.045 80.000 73.945 ;
        RECT 0.000 71.945 2.100 72.045 ;
        RECT 77.900 71.945 80.000 72.045 ;
        RECT 0.000 70.045 2.985 71.945 ;
        RECT 77.015 70.045 80.000 71.945 ;
        RECT 0.000 69.945 2.100 70.045 ;
        RECT 77.900 69.945 80.000 70.045 ;
        RECT 0.000 68.045 2.985 69.945 ;
        RECT 77.015 68.045 80.000 69.945 ;
        RECT 0.000 67.945 2.100 68.045 ;
        RECT 77.900 67.945 80.000 68.045 ;
        RECT 0.000 66.045 2.985 67.945 ;
        RECT 77.015 66.045 80.000 67.945 ;
        RECT 0.000 65.945 2.100 66.045 ;
        RECT 77.900 65.945 80.000 66.045 ;
        RECT 0.000 64.045 2.985 65.945 ;
        RECT 77.015 64.045 80.000 65.945 ;
        RECT 0.000 63.945 2.100 64.045 ;
        RECT 77.900 63.945 80.000 64.045 ;
        RECT 0.000 62.045 2.985 63.945 ;
        RECT 77.015 62.045 80.000 63.945 ;
        RECT 0.000 61.945 2.100 62.045 ;
        RECT 77.900 61.945 80.000 62.045 ;
        RECT 0.000 60.045 2.985 61.945 ;
        RECT 77.015 60.045 80.000 61.945 ;
        RECT 0.000 59.945 2.100 60.045 ;
        RECT 77.900 59.945 80.000 60.045 ;
        RECT 0.000 58.045 2.985 59.945 ;
        RECT 77.015 58.045 80.000 59.945 ;
        RECT 0.000 57.945 2.100 58.045 ;
        RECT 77.900 57.945 80.000 58.045 ;
        RECT 0.000 56.045 2.985 57.945 ;
        RECT 77.015 56.045 80.000 57.945 ;
        RECT 0.000 55.945 2.100 56.045 ;
        RECT 77.900 55.945 80.000 56.045 ;
        RECT 0.000 54.045 2.985 55.945 ;
        RECT 77.015 54.045 80.000 55.945 ;
        RECT 0.000 53.945 2.100 54.045 ;
        RECT 77.900 53.945 80.000 54.045 ;
        RECT 0.000 52.045 2.985 53.945 ;
        RECT 77.015 52.045 80.000 53.945 ;
        RECT 0.000 51.945 2.100 52.045 ;
        RECT 77.900 51.945 80.000 52.045 ;
        RECT 0.000 50.045 2.985 51.945 ;
        RECT 77.015 50.045 80.000 51.945 ;
        RECT 0.000 49.945 2.100 50.045 ;
        RECT 77.900 49.945 80.000 50.045 ;
        RECT 0.000 48.045 2.985 49.945 ;
        RECT 77.015 48.045 80.000 49.945 ;
        RECT 0.000 47.950 2.100 48.045 ;
        RECT 77.900 47.950 80.000 48.045 ;
        RECT 0.000 46.050 2.985 47.950 ;
        RECT 77.015 46.050 80.000 47.950 ;
        RECT 0.000 45.950 2.100 46.050 ;
        RECT 77.900 45.950 80.000 46.050 ;
        RECT 0.000 44.050 2.985 45.950 ;
        RECT 77.015 44.050 80.000 45.950 ;
        RECT 0.000 43.950 2.100 44.050 ;
        RECT 77.900 43.950 80.000 44.050 ;
        RECT 0.000 42.050 2.985 43.950 ;
        RECT 77.015 42.050 80.000 43.950 ;
        RECT 0.000 41.950 2.100 42.050 ;
        RECT 77.900 41.950 80.000 42.050 ;
        RECT 0.000 40.050 2.985 41.950 ;
        RECT 77.015 40.050 80.000 41.950 ;
        RECT 0.000 39.950 2.100 40.050 ;
        RECT 77.900 39.950 80.000 40.050 ;
        RECT 0.000 38.050 2.985 39.950 ;
        RECT 77.015 38.050 80.000 39.950 ;
        RECT 0.000 37.950 2.100 38.050 ;
        RECT 77.900 37.950 80.000 38.050 ;
        RECT 0.000 36.050 2.985 37.950 ;
        RECT 77.015 36.050 80.000 37.950 ;
        RECT 0.000 35.950 2.100 36.050 ;
        RECT 77.900 35.950 80.000 36.050 ;
        RECT 0.000 34.050 2.985 35.950 ;
        RECT 77.015 34.050 80.000 35.950 ;
        RECT 0.000 33.950 2.100 34.050 ;
        RECT 77.900 33.950 80.000 34.050 ;
        RECT 0.000 32.050 2.985 33.950 ;
        RECT 77.015 32.050 80.000 33.950 ;
        RECT 0.000 31.950 2.100 32.050 ;
        RECT 77.900 31.950 80.000 32.050 ;
        RECT 0.000 30.050 2.985 31.950 ;
        RECT 77.015 30.050 80.000 31.950 ;
        RECT 0.000 29.950 2.100 30.050 ;
        RECT 77.900 29.950 80.000 30.050 ;
        RECT 0.000 28.050 2.985 29.950 ;
        RECT 77.015 28.050 80.000 29.950 ;
        RECT 0.000 27.950 2.100 28.050 ;
        RECT 77.900 27.950 80.000 28.050 ;
        RECT 0.000 26.050 2.985 27.950 ;
        RECT 77.015 26.050 80.000 27.950 ;
        RECT 0.000 25.950 2.100 26.050 ;
        RECT 77.900 25.950 80.000 26.050 ;
        RECT 0.000 24.050 2.985 25.950 ;
        RECT 77.015 24.050 80.000 25.950 ;
        RECT 0.000 23.950 2.100 24.050 ;
        RECT 77.900 23.950 80.000 24.050 ;
        RECT 0.000 22.050 2.985 23.950 ;
        RECT 77.015 22.050 80.000 23.950 ;
        RECT 0.000 21.950 2.100 22.050 ;
        RECT 77.900 21.950 80.000 22.050 ;
        RECT 0.000 20.050 2.985 21.950 ;
        RECT 77.015 20.050 80.000 21.950 ;
        RECT 0.000 19.950 2.100 20.050 ;
        RECT 77.900 19.950 80.000 20.050 ;
        RECT 0.000 18.050 2.985 19.950 ;
        RECT 77.015 18.050 80.000 19.950 ;
        RECT 0.000 17.950 2.100 18.050 ;
        RECT 77.900 17.950 80.000 18.050 ;
        RECT 0.000 16.050 2.985 17.950 ;
        RECT 77.015 16.050 80.000 17.950 ;
        RECT 0.000 15.950 2.100 16.050 ;
        RECT 77.900 15.950 80.000 16.050 ;
        RECT 0.000 14.050 2.985 15.950 ;
        RECT 77.015 14.050 80.000 15.950 ;
        RECT 0.000 13.950 2.100 14.050 ;
        RECT 77.900 13.950 80.000 14.050 ;
        RECT 0.000 12.050 2.985 13.950 ;
        RECT 77.015 12.050 80.000 13.950 ;
        RECT 0.000 11.955 2.100 12.050 ;
        RECT 77.900 11.955 80.000 12.050 ;
        RECT 0.000 10.055 2.985 11.955 ;
        RECT 77.015 10.055 80.000 11.955 ;
        RECT 0.000 9.985 2.100 10.055 ;
        RECT 77.900 9.985 80.000 10.055 ;
        RECT 0.000 9.100 2.985 9.985 ;
        RECT 3.080 9.100 4.980 9.985 ;
        RECT 5.080 9.100 6.980 9.985 ;
        RECT 7.075 9.100 8.975 9.985 ;
        RECT 9.075 9.100 10.975 9.985 ;
        RECT 11.075 9.100 12.975 9.985 ;
        RECT 13.070 9.100 14.970 9.985 ;
        RECT 15.070 9.100 16.970 9.985 ;
        RECT 17.070 9.100 18.970 9.985 ;
        RECT 19.065 9.100 20.965 9.985 ;
        RECT 21.065 9.100 22.965 9.985 ;
        RECT 23.060 9.100 24.960 9.985 ;
        RECT 25.060 9.100 26.960 9.985 ;
        RECT 27.060 9.100 28.960 9.985 ;
        RECT 29.055 9.100 30.955 9.985 ;
        RECT 31.055 9.100 32.955 9.985 ;
        RECT 33.055 9.100 34.955 9.985 ;
        RECT 35.050 9.100 36.950 9.985 ;
        RECT 37.050 9.100 38.950 9.985 ;
        RECT 39.050 9.100 40.950 9.985 ;
        RECT 41.045 9.100 42.945 9.985 ;
        RECT 43.045 9.100 44.945 9.985 ;
        RECT 45.040 9.100 46.940 9.985 ;
        RECT 47.040 9.100 48.940 9.985 ;
        RECT 49.040 9.100 50.940 9.985 ;
        RECT 51.035 9.100 52.935 9.985 ;
        RECT 53.035 9.100 54.935 9.985 ;
        RECT 55.035 9.100 56.935 9.985 ;
        RECT 57.030 9.100 58.930 9.985 ;
        RECT 59.030 9.100 60.930 9.985 ;
        RECT 61.025 9.100 62.925 9.985 ;
        RECT 63.025 9.100 64.925 9.985 ;
        RECT 65.025 9.100 66.925 9.985 ;
        RECT 67.020 9.100 68.920 9.985 ;
        RECT 69.020 9.100 70.920 9.985 ;
        RECT 71.020 9.100 72.920 9.985 ;
        RECT 73.015 9.100 74.915 9.985 ;
        RECT 75.015 9.100 76.915 9.985 ;
        RECT 77.015 9.100 80.000 9.985 ;
        RECT 0.000 7.000 80.000 9.100 ;
        RECT 16.500 0.000 23.500 7.000 ;
        RECT 26.500 0.000 33.500 7.000 ;
        RECT 36.500 0.000 43.500 7.000 ;
        RECT 46.500 0.000 53.500 7.000 ;
        RECT 56.500 0.000 63.500 7.000 ;
  END
END sg13g2_bpd80

END LIBRARY
