VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.34 BY 6.12 ;
END obssite

#--------EOF---------

MACRO AN2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1
MACRO AN2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 1.390 0.815 2.210 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.210 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 0.335 2.690 ;
        RECT 0.175 2.530 2.735 2.690 ;
        RECT 2.525 2.530 2.785 2.690 ;
  END
END AN2D1_1
MACRO AN2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1_2
MACRO AN2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 2.255 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1_3
#--------EOF---------

MACRO AN2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1
MACRO AN2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 1.390 0.815 2.210 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.210 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 0.335 2.690 ;
        RECT 0.175 2.530 2.735 2.690 ;
        RECT 2.525 2.530 2.785 2.690 ;
  END
END AN2D1_1
MACRO AN2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1_2
MACRO AN2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 2.255 1.150 ;
        RECT 2.095 0.990 2.255 3.650 ;
        RECT 2.045 3.490 2.305 3.650 ;
  END
END AN2D1_3
#--------EOF---------

MACRO AO21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 1.775 3.650 ;
        RECT 1.565 3.490 1.825 3.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 2.575 2.530 2.735 3.650 ;
        RECT 2.525 3.490 2.785 3.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 1.295 1.150 ;
        RECT 1.135 0.990 1.295 3.170 ;
        RECT 1.085 3.010 1.345 3.170 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 3.055 0.990 3.215 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.170 0.335 4.790 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END AO21D1
MACRO AO21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.525 4.630 2.785 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 2.575 0.990 3.215 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 3.055 4.170 3.215 4.790 ;
  END
END AO21D1_1
MACRO AO21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 1.135 0.330 4.655 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AO21D1_2
MACRO AO21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
  END
END AO21D1_3
#--------EOF---------

MACRO AO21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 1.775 3.650 ;
        RECT 1.565 3.490 1.825 3.650 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 2.575 2.530 2.735 3.650 ;
        RECT 2.525 3.490 2.785 3.650 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 1.295 1.150 ;
        RECT 1.135 0.990 1.295 3.170 ;
        RECT 1.085 3.010 1.345 3.170 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 3.055 0.990 3.215 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.170 0.335 4.790 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END AO21D1
MACRO AO21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.525 4.630 2.785 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 2.575 0.990 3.215 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 3.055 4.170 3.215 4.790 ;
  END
END AO21D1_1
MACRO AO21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 1.135 0.330 4.655 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AO21D1_2
MACRO AO21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
  END
END AO21D1_3
#--------EOF---------

MACRO AOI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
  END
END AOI21D1
MACRO AOI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 4.630 3.215 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.630 1.295 5.130 ;
  END
END AOI21D1_1
MACRO AOI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 2.050 0.385 2.210 ;
        RECT 0.175 2.050 0.335 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.655 0.990 2.255 1.150 ;
        RECT 0.655 0.990 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 0.655 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AOI21D1_2
MACRO AOI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 0.175 4.170 0.335 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AOI21D1_3
#--------EOF---------

MACRO AOI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 2.255 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
  END
END AOI21D1
MACRO AOI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 4.630 3.215 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 1.135 4.630 1.295 5.130 ;
  END
END AOI21D1_1
MACRO AOI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 2.050 0.385 2.210 ;
        RECT 0.175 2.050 0.335 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.655 0.990 2.255 1.150 ;
        RECT 0.655 0.990 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 0.655 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AOI21D1_2
MACRO AOI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.170 2.255 4.330 ;
        RECT 0.175 4.170 0.335 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 4.630 1.295 5.130 ;
        RECT 1.135 4.970 3.215 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
  END
END AOI21D1_3
#--------EOF---------

MACRO BUFFD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 1.775 3.650 ;
        RECT 1.615 3.490 1.775 5.130 ;
        RECT 1.615 4.970 2.255 5.130 ;
        RECT 0.655 0.990 2.255 1.150 ;
        RECT 0.655 0.990 0.815 2.210 ;
        RECT 0.605 2.050 0.865 2.210 ;
  END
END BUFFD1
MACRO BUFFD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 0.655 3.490 1.775 3.650 ;
        RECT 0.655 3.490 0.815 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.990 1.775 2.210 ;
        RECT 1.565 2.050 1.825 2.210 ;
  END
END BUFFD1_1
#--------EOF---------

MACRO BUFFD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 1.775 3.650 ;
        RECT 1.615 3.490 1.775 5.130 ;
        RECT 1.615 4.970 2.255 5.130 ;
        RECT 0.655 0.990 2.255 1.150 ;
        RECT 0.655 0.990 0.815 2.210 ;
        RECT 0.605 2.050 0.865 2.210 ;
  END
END BUFFD1
MACRO BUFFD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 0.655 3.490 1.775 3.650 ;
        RECT 0.655 3.490 0.815 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.990 1.775 2.210 ;
        RECT 1.565 2.050 1.825 2.210 ;
  END
END BUFFD1_1
#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFCNQD1 0 0 ; 
  SIZE 17.000 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cdn
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 7.375 2.050 8.015 2.210 ;
    END 
  END cdn
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 16.445 0.990 16.705 1.150 ;
        RECT 15.485 4.630 15.745 4.790 ;
        RECT 16.495 0.990 16.655 4.330 ;
        RECT 15.535 4.170 16.655 4.330 ;
        RECT 15.535 4.170 15.695 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 8.815 4.970 8.975 6.050 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 12.655 4.970 12.815 6.050 ;
        RECT 0.000 5.970 17.000 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.855 0.070 8.015 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.655 0.070 12.815 1.150 ;
        RECT 15.485 0.990 15.745 1.150 ;
        RECT 15.535 0.070 15.695 1.150 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.330 1.775 1.150 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 10.415 3.170 ;
        RECT 10.205 3.010 10.465 3.170 ;
        RECT 0.175 4.970 0.335 5.790 ;
        RECT 0.175 5.630 1.775 5.790 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 5.130 ;
        RECT 2.045 4.170 2.305 4.330 ;
        RECT 2.095 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 3.535 3.490 5.615 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 8.765 3.490 9.025 3.650 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 2.690 ;
        RECT 4.975 2.530 9.455 2.690 ;
        RECT 9.245 2.530 9.505 2.690 ;
        RECT 8.285 2.530 8.545 2.690 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 4.975 4.170 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 4.925 2.530 5.185 2.690 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 5.935 4.970 8.015 5.130 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 8.815 0.990 8.975 1.550 ;
        RECT 6.415 1.390 8.975 1.550 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.365 4.170 6.625 4.330 ;
        RECT 6.415 4.170 9.935 4.330 ;
        RECT 9.775 4.170 9.935 4.790 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 10.685 4.630 10.945 4.790 ;
        RECT 9.775 0.330 9.935 1.150 ;
        RECT 9.775 0.330 12.335 0.490 ;
        RECT 12.125 0.330 12.385 0.490 ;
        RECT 14.045 2.050 14.305 2.210 ;
        RECT 14.095 2.050 14.255 4.330 ;
        RECT 10.735 4.170 14.255 4.330 ;
        RECT 10.735 4.170 10.895 4.790 ;
        RECT 14.045 3.490 14.305 3.650 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.735 0.990 11.855 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 12.125 1.390 12.385 1.550 ;
        RECT 12.175 1.390 14.735 1.550 ;
        RECT 14.575 0.990 14.735 1.550 ;
        RECT 14.575 1.390 14.735 4.790 ;
        RECT 13.615 4.630 14.735 4.790 ;
  END
END DFCNQD1
#--------EOF---------

MACRO DFCNQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFCNQD1_1 0 0 ; 
  SIZE 17.000 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cdn
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 7.375 2.050 8.015 2.210 ;
    END 
  END cdn
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 16.445 0.990 16.705 1.150 ;
        RECT 15.485 4.630 15.745 4.790 ;
        RECT 16.495 0.990 16.655 4.330 ;
        RECT 15.535 4.170 16.655 4.330 ;
        RECT 15.535 4.170 15.695 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 8.765 4.970 9.025 5.130 ;
        RECT 8.815 4.970 8.975 6.050 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 12.655 4.970 12.815 6.050 ;
        RECT 0.000 5.970 17.000 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.855 0.070 8.015 1.150 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.655 0.070 12.815 1.150 ;
        RECT 15.485 0.990 15.745 1.150 ;
        RECT 15.535 0.070 15.695 1.150 ;
        RECT 0.000 -0.150 17.000 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.330 1.775 1.150 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 10.415 3.170 ;
        RECT 10.205 3.010 10.465 3.170 ;
        RECT 0.175 4.970 0.335 5.790 ;
        RECT 0.175 5.630 1.775 5.790 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 5.130 ;
        RECT 2.045 4.170 2.305 4.330 ;
        RECT 2.095 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 3.535 3.490 5.615 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 8.765 3.490 9.025 3.650 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 2.690 ;
        RECT 4.975 2.530 9.455 2.690 ;
        RECT 9.245 2.530 9.505 2.690 ;
        RECT 8.285 2.530 8.545 2.690 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 4.975 4.170 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 4.925 2.530 5.185 2.690 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 7.805 4.970 8.065 5.130 ;
        RECT 5.935 4.970 8.015 5.130 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 8.815 0.990 8.975 1.550 ;
        RECT 6.415 1.390 8.975 1.550 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.365 4.170 6.625 4.330 ;
        RECT 6.415 4.170 9.935 4.330 ;
        RECT 9.775 4.170 9.935 4.790 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 10.685 4.630 10.945 4.790 ;
        RECT 9.775 0.330 9.935 1.150 ;
        RECT 9.775 0.330 12.335 0.490 ;
        RECT 12.125 0.330 12.385 0.490 ;
        RECT 14.045 2.050 14.305 2.210 ;
        RECT 14.095 2.050 14.255 4.330 ;
        RECT 10.735 4.170 14.255 4.330 ;
        RECT 10.735 4.170 10.895 4.790 ;
        RECT 14.045 3.490 14.305 3.650 ;
        RECT 10.685 0.990 10.945 1.150 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.735 0.990 11.855 1.150 ;
        RECT 14.525 0.990 14.785 1.150 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 12.125 1.390 12.385 1.550 ;
        RECT 12.175 1.390 14.735 1.550 ;
        RECT 14.575 0.990 14.735 1.550 ;
        RECT 14.575 1.390 14.735 4.790 ;
        RECT 13.615 4.630 14.735 4.790 ;
  END
END DFCNQD1_1
#--------EOF---------

MACRO DFQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1 0 0 ; 
  SIZE 14.960 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 0.655 2.530 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 13.615 0.990 13.775 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.960 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.960 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.125 3.010 0.385 3.170 ;
        RECT 0.175 3.010 0.335 4.790 ;
        RECT 12.125 0.330 12.385 0.490 ;
        RECT 7.855 0.330 12.335 0.490 ;
        RECT 7.805 0.330 8.065 0.490 ;
        RECT 0.175 0.990 0.335 3.170 ;
        RECT 0.175 3.010 0.335 4.330 ;
        RECT 0.175 4.170 3.215 4.330 ;
        RECT 3.005 4.170 3.265 4.330 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 4.015 3.490 5.615 3.650 ;
        RECT 4.015 3.490 4.175 4.330 ;
        RECT 3.965 4.170 4.225 4.330 ;
        RECT 5.405 5.630 5.665 5.790 ;
        RECT 3.535 5.630 5.615 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 10.735 0.990 12.815 1.150 ;
        RECT 10.735 0.990 10.895 1.550 ;
        RECT 6.895 1.390 10.895 1.550 ;
        RECT 6.895 0.990 7.055 1.550 ;
        RECT 9.295 1.390 9.455 3.650 ;
        RECT 9.245 3.490 9.505 3.650 ;
        RECT 9.245 2.050 9.505 2.210 ;
        RECT 9.295 2.050 9.455 4.790 ;
        RECT 9.295 4.630 12.815 4.790 ;
        RECT 12.655 4.630 12.815 5.130 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.055 2.050 8.495 2.210 ;
        RECT 8.285 2.050 8.545 2.210 ;
        RECT 8.285 3.010 8.545 3.170 ;
        RECT 3.535 3.010 8.495 3.170 ;
        RECT 3.535 3.010 3.695 4.790 ;
        RECT 3.055 4.630 3.695 4.790 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 3.485 1.390 3.745 1.550 ;
        RECT 3.535 1.390 6.095 1.550 ;
        RECT 5.935 0.990 6.095 1.550 ;
        RECT 6.365 4.630 6.625 4.790 ;
        RECT 5.935 4.630 6.575 4.790 ;
        RECT 5.935 1.390 6.575 1.550 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 4.630 6.575 5.790 ;
        RECT 6.415 5.630 12.335 5.790 ;
        RECT 12.125 5.630 12.385 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 7.535 0.490 ;
        RECT 7.375 0.330 7.535 1.150 ;
        RECT 7.375 0.990 8.015 1.150 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 4.495 4.170 8.015 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.165 1.390 11.425 1.550 ;
        RECT 11.215 1.390 13.295 1.550 ;
        RECT 13.085 1.390 13.345 1.550 ;
        RECT 10.205 0.990 10.465 1.150 ;
        RECT 9.775 0.990 10.415 1.150 ;
  END
END DFQD1
MACRO DFQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_1 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 0.175 0.330 1.775 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 9.245 2.050 9.505 2.210 ;
        RECT 9.295 2.050 9.455 3.650 ;
        RECT 9.245 3.490 9.505 3.650 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 0.335 5.790 ;
        RECT 0.175 5.630 3.695 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.775 3.490 9.935 4.330 ;
        RECT 8.815 4.170 9.935 4.330 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 3.055 2.530 7.535 2.690 ;
        RECT 7.325 2.530 7.585 2.690 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 3.055 2.050 7.535 2.210 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 3.485 4.170 3.745 4.330 ;
        RECT 3.535 4.170 3.695 4.790 ;
        RECT 3.535 4.630 6.095 4.790 ;
        RECT 8.285 0.330 8.545 0.490 ;
        RECT 5.935 0.330 8.495 0.490 ;
        RECT 5.935 0.330 6.095 1.150 ;
        RECT 5.935 4.630 6.095 5.790 ;
        RECT 5.935 5.630 9.455 5.790 ;
        RECT 9.245 5.630 9.505 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 4.495 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 7.855 1.390 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_1
MACRO DFQD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_2 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.990 1.775 2.210 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.295 3.490 9.935 3.650 ;
        RECT 9.295 3.490 9.455 4.790 ;
        RECT 8.815 4.630 9.455 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 4.975 0.330 7.535 0.490 ;
        RECT 7.325 0.330 7.585 0.490 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 4.975 4.170 7.535 4.330 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 5.405 1.390 5.665 1.550 ;
        RECT 2.095 1.390 5.615 1.550 ;
        RECT 2.095 0.990 2.255 1.550 ;
        RECT 8.285 2.050 8.545 2.210 ;
        RECT 2.575 2.050 8.495 2.210 ;
        RECT 2.575 2.050 2.735 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 5.455 1.390 5.615 2.210 ;
        RECT 8.335 2.050 8.495 5.790 ;
        RECT 8.335 5.630 9.455 5.790 ;
        RECT 9.245 5.630 9.505 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 3.535 5.630 8.495 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 6.365 3.490 6.625 3.650 ;
        RECT 6.415 3.490 8.015 3.650 ;
        RECT 7.855 3.490 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_2
MACRO DFQD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_3 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 3.010 1.345 3.170 ;
        RECT 1.135 3.010 1.295 3.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 9.245 0.330 9.505 0.490 ;
        RECT 4.015 0.330 9.455 0.490 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 2.575 0.990 4.175 1.150 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 1.775 2.210 ;
        RECT 1.615 2.050 1.775 4.790 ;
        RECT 1.615 4.630 2.255 4.790 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 0.655 2.530 2.255 2.690 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.295 3.490 9.935 3.650 ;
        RECT 9.295 3.490 9.455 4.790 ;
        RECT 8.815 4.630 9.455 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 4.975 2.050 7.535 2.210 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.175 0.330 3.695 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 8.495 5.130 ;
        RECT 8.335 3.490 8.495 5.130 ;
        RECT 8.285 3.490 8.545 3.650 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 3.535 4.970 3.695 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 7.855 1.390 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_3
#--------EOF---------

MACRO DFQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1 0 0 ; 
  SIZE 14.960 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 0.655 2.530 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 13.565 0.990 13.825 1.150 ;
        RECT 13.565 4.630 13.825 4.790 ;
        RECT 13.615 0.990 13.775 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.960 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.960 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.125 3.010 0.385 3.170 ;
        RECT 0.175 3.010 0.335 4.790 ;
        RECT 12.125 0.330 12.385 0.490 ;
        RECT 7.855 0.330 12.335 0.490 ;
        RECT 7.805 0.330 8.065 0.490 ;
        RECT 0.175 0.990 0.335 3.170 ;
        RECT 0.175 3.010 0.335 4.330 ;
        RECT 0.175 4.170 3.215 4.330 ;
        RECT 3.005 4.170 3.265 4.330 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 4.015 3.490 5.615 3.650 ;
        RECT 4.015 3.490 4.175 4.330 ;
        RECT 3.965 4.170 4.225 4.330 ;
        RECT 5.405 5.630 5.665 5.790 ;
        RECT 3.535 5.630 5.615 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 12.605 4.970 12.865 5.130 ;
        RECT 10.735 0.990 12.815 1.150 ;
        RECT 10.735 0.990 10.895 1.550 ;
        RECT 6.895 1.390 10.895 1.550 ;
        RECT 6.895 0.990 7.055 1.550 ;
        RECT 9.295 1.390 9.455 3.650 ;
        RECT 9.245 3.490 9.505 3.650 ;
        RECT 9.245 2.050 9.505 2.210 ;
        RECT 9.295 2.050 9.455 4.790 ;
        RECT 9.295 4.630 12.815 4.790 ;
        RECT 12.655 4.630 12.815 5.130 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.055 2.050 8.495 2.210 ;
        RECT 8.285 2.050 8.545 2.210 ;
        RECT 8.285 3.010 8.545 3.170 ;
        RECT 3.535 3.010 8.495 3.170 ;
        RECT 3.535 3.010 3.695 4.790 ;
        RECT 3.055 4.630 3.695 4.790 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 3.485 1.390 3.745 1.550 ;
        RECT 3.535 1.390 6.095 1.550 ;
        RECT 5.935 0.990 6.095 1.550 ;
        RECT 6.365 4.630 6.625 4.790 ;
        RECT 5.935 4.630 6.575 4.790 ;
        RECT 5.935 1.390 6.575 1.550 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 4.630 6.575 5.790 ;
        RECT 6.415 5.630 12.335 5.790 ;
        RECT 12.125 5.630 12.385 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 7.535 0.490 ;
        RECT 7.375 0.330 7.535 1.150 ;
        RECT 7.375 0.990 8.015 1.150 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 4.495 4.170 8.015 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
        RECT 9.725 0.990 9.985 1.150 ;
        RECT 11.165 1.390 11.425 1.550 ;
        RECT 11.215 1.390 13.295 1.550 ;
        RECT 13.085 1.390 13.345 1.550 ;
        RECT 10.205 0.990 10.465 1.150 ;
        RECT 9.775 0.990 10.415 1.150 ;
  END
END DFQD1
MACRO DFQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_1 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 0.175 0.330 1.775 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 9.245 2.050 9.505 2.210 ;
        RECT 9.295 2.050 9.455 3.650 ;
        RECT 9.245 3.490 9.505 3.650 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 0.335 5.790 ;
        RECT 0.175 5.630 3.695 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.775 3.490 9.935 4.330 ;
        RECT 8.815 4.170 9.935 4.330 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 3.055 2.530 7.535 2.690 ;
        RECT 7.325 2.530 7.585 2.690 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 3.055 2.050 7.535 2.210 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 3.485 4.170 3.745 4.330 ;
        RECT 3.535 4.170 3.695 4.790 ;
        RECT 3.535 4.630 6.095 4.790 ;
        RECT 8.285 0.330 8.545 0.490 ;
        RECT 5.935 0.330 8.495 0.490 ;
        RECT 5.935 0.330 6.095 1.150 ;
        RECT 5.935 4.630 6.095 5.790 ;
        RECT 5.935 5.630 9.455 5.790 ;
        RECT 9.245 5.630 9.505 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 4.495 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 7.855 1.390 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_1
MACRO DFQD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_2 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 1.775 1.150 ;
        RECT 1.615 0.990 1.775 2.210 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.295 3.490 9.935 3.650 ;
        RECT 9.295 3.490 9.455 4.790 ;
        RECT 8.815 4.630 9.455 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 4.975 0.330 7.535 0.490 ;
        RECT 7.325 0.330 7.585 0.490 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 4.975 4.170 7.535 4.330 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 5.405 1.390 5.665 1.550 ;
        RECT 2.095 1.390 5.615 1.550 ;
        RECT 2.095 0.990 2.255 1.550 ;
        RECT 8.285 2.050 8.545 2.210 ;
        RECT 2.575 2.050 8.495 2.210 ;
        RECT 2.575 2.050 2.735 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 5.455 1.390 5.615 2.210 ;
        RECT 8.335 2.050 8.495 5.790 ;
        RECT 8.335 5.630 9.455 5.790 ;
        RECT 9.245 5.630 9.505 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 3.535 5.630 8.495 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 6.365 3.490 6.625 3.650 ;
        RECT 6.415 3.490 8.015 3.650 ;
        RECT 7.855 3.490 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_2
MACRO DFQD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_3 0 0 ; 
  SIZE 14.280 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN cp
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 3.010 1.345 3.170 ;
        RECT 1.135 3.010 1.295 3.650 ;
    END 
  END cp
  PIN d
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END d
  PIN q
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 12.605 0.990 12.865 1.150 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 12.655 0.990 12.815 4.790 ;
    END 
  END q
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 14.280 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 14.280 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 9.245 0.330 9.505 0.490 ;
        RECT 4.015 0.330 9.455 0.490 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 2.575 0.990 4.175 1.150 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 1.775 2.210 ;
        RECT 1.615 2.050 1.775 4.790 ;
        RECT 1.615 4.630 2.255 4.790 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 0.655 2.530 2.255 2.690 ;
        RECT 0.605 2.530 0.865 2.690 ;
        RECT 8.765 0.990 9.025 1.150 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 8.815 0.990 11.375 1.150 ;
        RECT 11.215 0.330 11.375 1.150 ;
        RECT 11.165 0.330 11.425 0.490 ;
        RECT 9.775 0.990 9.935 3.650 ;
        RECT 9.775 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
        RECT 9.295 3.490 9.935 3.650 ;
        RECT 9.295 3.490 9.455 4.790 ;
        RECT 8.815 4.630 9.455 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
        RECT 7.325 2.050 7.585 2.210 ;
        RECT 4.975 2.050 7.535 2.210 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.175 0.330 3.695 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 8.495 5.130 ;
        RECT 8.335 3.490 8.495 5.130 ;
        RECT 8.285 3.490 8.545 3.650 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 3.535 4.970 3.695 5.790 ;
        RECT 7.805 0.990 8.065 1.150 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 6.365 1.390 6.625 1.550 ;
        RECT 6.415 1.390 8.015 1.550 ;
        RECT 7.855 0.990 8.015 1.550 ;
        RECT 7.855 1.390 8.015 4.790 ;
        RECT 11.645 0.990 11.905 1.150 ;
        RECT 10.205 1.390 10.465 1.550 ;
        RECT 10.255 1.390 12.335 1.550 ;
        RECT 12.175 0.330 12.335 1.550 ;
        RECT 12.175 0.330 13.295 0.490 ;
        RECT 13.085 0.330 13.345 0.490 ;
        RECT 11.695 0.990 11.855 1.550 ;
  END
END DFQD1_3
#--------EOF---------

MACRO FILL1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL1 0 0 ; 
  SIZE 0.340 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 0.340 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.340 0.150 ;
    END 
  END vss 
END FILL1
#--------EOF---------

MACRO FILL1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL1 0 0 ; 
  SIZE 0.340 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 0.340 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.340 0.150 ;
    END 
  END vss 
END FILL1
#--------EOF---------

MACRO FILL2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL2 0 0 ; 
  SIZE 0.680 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 0.680 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.680 0.150 ;
    END 
  END vss 
END FILL2
#--------EOF---------

MACRO FILL2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL2 0 0 ; 
  SIZE 0.680 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 0.680 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 0.680 0.150 ;
    END 
  END vss 
END FILL2
#--------EOF---------

MACRO FILL4
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL4 0 0 ; 
  SIZE 1.360 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 1.360 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 1.360 0.150 ;
    END 
  END vss 
END FILL4
#--------EOF---------

MACRO FILL4
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL4 0 0 ; 
  SIZE 1.360 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 1.360 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 1.360 0.150 ;
    END 
  END vss 
END FILL4
#--------EOF---------

MACRO FILL8
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL8 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END FILL8
#--------EOF---------

MACRO FILL8
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL8 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END FILL8
#--------EOF---------

MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1
MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1
MACRO INVD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_1
MACRO INVD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_2 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_2
MACRO INVD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_3 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_3
#--------EOF---------

MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1
MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1
MACRO INVD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_1 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_1
MACRO INVD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_2 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_2
MACRO INVD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1_3 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
END INVD1_3
#--------EOF---------

MACRO MUX2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 1.390 2.735 2.210 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.210 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 0.655 0.330 4.655 0.490 ;
        RECT 4.495 0.330 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 5.405 2.050 5.665 2.210 ;
        RECT 5.455 2.050 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 2.210 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 1.135 3.490 1.295 4.790 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.015 0.990 4.175 3.650 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 0.175 2.530 2.735 2.690 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 4.015 2.530 4.175 5.130 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.925 0.330 5.185 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 3.005 5.630 3.265 5.790 ;
        RECT 3.055 5.630 5.135 5.790 ;
        RECT 4.975 4.970 5.135 5.790 ;
  END
END MUX2D1
MACRO MUX2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 3.055 3.010 4.655 3.170 ;
        RECT 3.005 3.010 3.265 3.170 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 2.095 4.970 4.655 5.130 ;
        RECT 4.495 4.170 4.655 5.130 ;
        RECT 4.495 4.170 5.135 4.330 ;
        RECT 4.925 4.170 5.185 4.330 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.690 ;
        RECT 2.575 2.530 3.215 2.690 ;
        RECT 2.575 2.530 2.735 4.790 ;
        RECT 2.575 4.630 3.215 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 1.615 2.050 2.735 2.210 ;
        RECT 1.615 2.050 1.775 3.650 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 4.975 0.990 5.615 1.150 ;
        RECT 5.455 0.990 5.615 5.130 ;
        RECT 4.975 4.970 5.615 5.130 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 1.615 5.630 5.135 5.790 ;
        RECT 4.975 4.970 5.135 5.790 ;
  END
END MUX2D1_1
MACRO MUX2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.935 0.070 6.095 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 3.215 4.790 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 4.015 0.330 5.135 0.490 ;
        RECT 4.925 0.330 5.185 0.490 ;
        RECT 4.015 0.990 4.175 5.130 ;
        RECT 0.655 3.010 4.175 3.170 ;
        RECT 0.655 3.010 0.815 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
        RECT 0.175 0.990 0.335 3.170 ;
        RECT 0.175 3.010 0.815 3.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 2.210 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 1.135 3.490 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.445 0.990 4.705 1.150 ;
        RECT 4.495 0.990 5.135 1.150 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 3.535 0.330 3.695 2.690 ;
        RECT 3.485 2.530 3.745 2.690 ;
        RECT 4.975 0.990 5.135 5.130 ;
  END
END MUX2D1_2
MACRO MUX2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 2.735 1.150 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 4.970 4.175 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 3.215 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 5.130 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 2.095 3.010 4.655 3.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 2.575 4.170 2.735 5.130 ;
        RECT 2.575 4.970 3.695 5.130 ;
        RECT 3.535 4.630 3.695 5.130 ;
        RECT 3.535 4.630 5.135 4.790 ;
        RECT 4.975 4.630 5.135 5.130 ;
        RECT 4.975 0.990 5.135 4.790 ;
  END
END MUX2D1_3
#--------EOF---------

MACRO MUX2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 1.390 2.735 2.210 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 1.390 1.775 2.210 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 0.655 0.330 4.655 0.490 ;
        RECT 4.495 0.330 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 5.405 2.050 5.665 2.210 ;
        RECT 5.455 2.050 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 2.210 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 1.135 3.490 1.295 4.790 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.015 0.990 4.175 3.650 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 0.175 2.530 2.735 2.690 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 4.015 2.530 4.175 5.130 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.925 0.330 5.185 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 3.005 5.630 3.265 5.790 ;
        RECT 3.055 5.630 5.135 5.790 ;
        RECT 4.975 4.970 5.135 5.790 ;
  END
END MUX2D1
MACRO MUX2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 3.055 3.010 4.655 3.170 ;
        RECT 3.005 3.010 3.265 3.170 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 2.095 4.970 4.655 5.130 ;
        RECT 4.495 4.170 4.655 5.130 ;
        RECT 4.495 4.170 5.135 4.330 ;
        RECT 4.925 4.170 5.185 4.330 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.690 ;
        RECT 2.575 2.530 3.215 2.690 ;
        RECT 2.575 2.530 2.735 4.790 ;
        RECT 2.575 4.630 3.215 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 1.615 2.050 2.735 2.210 ;
        RECT 1.615 2.050 1.775 3.650 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 4.975 0.990 5.615 1.150 ;
        RECT 5.455 0.990 5.615 5.130 ;
        RECT 4.975 4.970 5.615 5.130 ;
        RECT 1.565 5.630 1.825 5.790 ;
        RECT 1.615 5.630 5.135 5.790 ;
        RECT 4.975 4.970 5.135 5.790 ;
  END
END MUX2D1_1
MACRO MUX2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.935 0.070 6.095 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 3.215 4.790 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 4.015 0.330 5.135 0.490 ;
        RECT 4.925 0.330 5.185 0.490 ;
        RECT 4.015 0.990 4.175 5.130 ;
        RECT 0.655 3.010 4.175 3.170 ;
        RECT 0.655 3.010 0.815 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
        RECT 0.175 0.990 0.335 3.170 ;
        RECT 0.175 3.010 0.815 3.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 2.210 ;
        RECT 1.085 2.050 1.345 2.210 ;
        RECT 1.085 3.490 1.345 3.650 ;
        RECT 1.135 3.490 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.445 0.990 4.705 1.150 ;
        RECT 4.495 0.990 5.135 1.150 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 3.535 0.330 3.695 2.690 ;
        RECT 3.485 2.530 3.745 2.690 ;
        RECT 4.975 0.990 5.135 5.130 ;
  END
END MUX2D1_2
MACRO MUX2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN i0
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END i0
  PIN i1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END i1
  PIN s
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 2.735 1.150 ;
    END 
  END s
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 4.970 4.175 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 3.215 4.790 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 5.130 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 2.095 3.010 4.655 3.170 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 2.575 4.170 2.735 5.130 ;
        RECT 2.575 4.970 3.695 5.130 ;
        RECT 3.535 4.630 3.695 5.130 ;
        RECT 3.535 4.630 5.135 4.790 ;
        RECT 4.975 4.630 5.135 5.130 ;
        RECT 4.975 0.990 5.135 4.790 ;
  END
END MUX2D1_3
#--------EOF---------

MACRO ND2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 1.135 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1
MACRO ND2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_1
MACRO ND2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_2
MACRO ND2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_3
#--------EOF---------

MACRO ND2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 1.135 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1
MACRO ND2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_1
MACRO ND2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_2
MACRO ND2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END ND2D1_3
#--------EOF---------

MACRO ND3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END ND3D1
MACRO ND3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_1 0 0 ; 
  SIZE 3.400 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.400 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.400 0.150 ;
    END 
  END vss 
END ND3D1_1
MACRO ND3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_2 0 0 ; 
  SIZE 4.760 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 0.175 0.330 4.175 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END ND3D1_2
MACRO ND3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END ND3D1_3
#--------EOF---------

MACRO ND3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END ND3D1
MACRO ND3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_1 0 0 ; 
  SIZE 3.400 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.400 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.400 0.150 ;
    END 
  END vss 
END ND3D1_1
MACRO ND3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_2 0 0 ; 
  SIZE 4.760 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.760 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.760 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 0.175 0.330 4.175 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END ND3D1_2
MACRO ND3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END ND3D1_3
#--------EOF---------

MACRO ND4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 0.990 3.215 4.330 ;
        RECT 3.055 4.170 4.175 4.330 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 0.175 0.330 4.175 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END ND4D1
MACRO ND4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.535 4.630 4.175 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 5.135 6.050 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 5.135 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
  END
END ND4D1_1
MACRO ND4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
END ND4D1_2
MACRO ND4D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 4.975 0.990 5.135 4.330 ;
        RECT 4.015 4.170 5.135 4.330 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 5.135 6.050 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 3.215 1.150 ;
  END
END ND4D1_3
#--------EOF---------

MACRO ND4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.055 0.990 3.215 4.330 ;
        RECT 3.055 4.170 4.175 4.330 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 1.135 4.170 3.215 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 0.175 0.330 4.175 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END ND4D1
MACRO ND4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.535 4.630 4.175 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 5.135 6.050 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 0.175 0.330 5.135 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
  END
END ND4D1_1
MACRO ND4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
END ND4D1_2
MACRO ND4D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 4.975 0.990 5.135 4.330 ;
        RECT 4.015 4.170 5.135 4.330 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 1.135 4.170 4.175 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 5.135 6.050 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 3.215 1.150 ;
  END
END ND4D1_3
#--------EOF---------

MACRO NR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 0.175 4.630 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1
MACRO NR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_1
MACRO NR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_2
MACRO NR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_3
#--------EOF---------

MACRO NR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 0.175 4.630 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 4.630 2.255 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1
MACRO NR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_1 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.095 0.070 2.255 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_1
MACRO NR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_2 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_2
MACRO NR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_3 0 0 ; 
  SIZE 2.720 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 2.720 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 2.720 0.150 ;
    END 
  END vss 
END NR2D1_3
#--------EOF---------

MACRO NR3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 1.615 0.330 1.775 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 2.735 1.150 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 3.055 0.990 3.215 3.650 ;
        RECT 1.135 3.490 3.215 3.650 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 0.175 4.970 8.015 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
  END
END NR3D1
MACRO NR3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_1 0 0 ; 
  SIZE 10.540 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 1.390 3.695 2.210 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 5.615 2.690 ;
        RECT 5.405 2.530 5.665 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 10.540 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 10.540 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 8.815 4.630 8.975 5.130 ;
        RECT 2.095 4.970 8.975 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 9.775 4.170 9.935 4.790 ;
        RECT 6.895 4.170 9.935 4.330 ;
        RECT 6.895 4.170 7.055 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 4.630 5.135 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
        RECT 1.615 4.170 3.215 4.330 ;
        RECT 1.615 4.170 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR3D1_1
MACRO NR3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_2 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 0.335 4.330 ;
        RECT 0.175 4.170 1.295 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 0.175 4.970 8.015 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
  END
END NR3D1_2
MACRO NR3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_3 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 1.135 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 3.055 4.970 8.015 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 2.575 4.170 4.175 4.330 ;
        RECT 2.575 4.170 2.735 5.130 ;
        RECT 0.175 4.970 2.735 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR3D1_3
#--------EOF---------

MACRO NR3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 1.615 0.330 1.775 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 2.735 1.150 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 3.055 0.990 3.215 3.650 ;
        RECT 1.135 3.490 3.215 3.650 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 0.175 4.970 8.015 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
  END
END NR3D1
MACRO NR3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_1 0 0 ; 
  SIZE 10.540 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 1.390 3.695 2.210 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 5.615 2.690 ;
        RECT 5.405 2.530 5.665 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 0.990 3.215 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 10.540 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 10.540 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 8.815 4.630 8.975 5.130 ;
        RECT 2.095 4.970 8.975 5.130 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 9.775 4.170 9.935 4.790 ;
        RECT 6.895 4.170 9.935 4.330 ;
        RECT 6.895 4.170 7.055 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 4.630 5.135 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.055 4.170 3.215 4.790 ;
        RECT 1.615 4.170 3.215 4.330 ;
        RECT 1.615 4.170 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR3D1_1
MACRO NR3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_2 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 0.175 0.990 0.335 4.330 ;
        RECT 0.175 4.170 1.295 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 0.175 4.970 8.015 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 4.175 4.790 ;
  END
END NR3D1_2
MACRO NR3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_3 0 0 ; 
  SIZE 9.520 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a3
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 3.215 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 1.135 0.990 2.255 1.150 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 9.520 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 9.520 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 7.855 4.630 8.015 5.130 ;
        RECT 3.055 4.970 8.015 5.130 ;
        RECT 3.055 4.630 3.215 5.130 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 8.815 4.170 8.975 4.790 ;
        RECT 5.935 4.170 8.975 4.330 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 2.575 4.170 4.175 4.330 ;
        RECT 2.575 4.170 2.735 5.130 ;
        RECT 0.175 4.970 2.735 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR3D1_3
#--------EOF---------

MACRO NR4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 0.655 0.330 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 4.015 3.490 6.575 3.650 ;
        RECT 6.365 3.490 6.625 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.490 8.065 3.650 ;
        RECT 7.855 3.490 12.335 3.650 ;
        RECT 12.125 3.490 12.385 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 4.630 11.855 4.790 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 12.175 4.630 12.815 4.790 ;
        RECT 12.175 4.170 12.335 4.790 ;
        RECT 7.855 4.170 12.335 4.330 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.630 3.215 4.790 ;
        RECT 1.615 4.630 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 4.975 4.630 6.575 4.790 ;
        RECT 6.415 4.170 6.575 4.790 ;
        RECT 6.415 4.170 7.535 4.330 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 7.325 4.970 7.585 5.130 ;
        RECT 7.375 4.970 9.935 5.130 ;
        RECT 9.775 4.630 9.935 5.130 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 2.095 4.170 6.095 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END NR4D1
MACRO NR4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_1 0 0 ; 
  SIZE 12.240 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 5.615 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 3.490 7.105 3.650 ;
        RECT 6.895 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 3.215 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 10.685 4.630 10.945 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 4.630 10.895 4.790 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 11.215 4.630 11.855 4.790 ;
        RECT 11.215 4.170 11.375 4.790 ;
        RECT 6.895 4.170 11.375 4.330 ;
        RECT 6.895 4.170 7.055 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 4.015 4.630 5.615 4.790 ;
        RECT 5.455 4.170 5.615 4.790 ;
        RECT 5.455 4.170 6.575 4.330 ;
        RECT 6.365 4.170 6.625 4.330 ;
        RECT 6.365 4.970 6.625 5.130 ;
        RECT 6.415 4.970 8.975 5.130 ;
        RECT 8.815 4.630 8.975 5.130 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 1.615 4.170 5.135 4.330 ;
        RECT 1.615 4.170 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR4D1_1
MACRO NR4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_2 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 4.655 5.790 ;
        RECT 3.535 5.630 4.655 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 4.445 5.630 4.705 5.790 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.655 0.330 3.695 0.490 ;
        RECT 0.655 0.330 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 3.695 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.490 8.065 3.650 ;
        RECT 7.855 3.490 12.335 3.650 ;
        RECT 12.125 3.490 12.385 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 4.630 11.855 4.790 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 12.175 4.630 12.815 4.790 ;
        RECT 12.175 4.170 12.335 4.790 ;
        RECT 7.855 4.170 12.335 4.330 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 4.630 3.215 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 2.095 4.170 2.735 4.330 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 7.325 4.970 7.585 5.130 ;
        RECT 7.375 4.970 9.935 5.130 ;
        RECT 9.775 4.630 9.935 5.130 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 6.095 4.790 ;
  END
END NR4D1_2
#--------EOF---------

MACRO NR4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 0.655 0.330 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 4.015 3.490 6.575 3.650 ;
        RECT 6.365 3.490 6.625 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.490 8.065 3.650 ;
        RECT 7.855 3.490 12.335 3.650 ;
        RECT 12.125 3.490 12.385 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 4.630 11.855 4.790 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 12.175 4.630 12.815 4.790 ;
        RECT 12.175 4.170 12.335 4.790 ;
        RECT 7.855 4.170 12.335 4.330 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 1.615 4.630 3.215 4.790 ;
        RECT 1.615 4.630 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 4.975 4.630 6.575 4.790 ;
        RECT 6.415 4.170 6.575 4.790 ;
        RECT 6.415 4.170 7.535 4.330 ;
        RECT 7.325 4.170 7.585 4.330 ;
        RECT 7.325 4.970 7.585 5.130 ;
        RECT 7.375 4.970 9.935 5.130 ;
        RECT 9.775 4.630 9.935 5.130 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 5.935 4.170 6.095 4.790 ;
        RECT 2.095 4.170 6.095 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END NR4D1
MACRO NR4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_1 0 0 ; 
  SIZE 12.240 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 3.490 3.265 3.650 ;
        RECT 3.055 3.490 5.615 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 3.490 7.105 3.650 ;
        RECT 6.895 3.490 11.375 3.650 ;
        RECT 11.165 3.490 11.425 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 3.215 1.150 ;
        RECT 1.135 0.990 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 12.240 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 12.240 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 10.685 4.630 10.945 4.790 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 4.630 10.895 4.790 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 11.215 4.630 11.855 4.790 ;
        RECT 11.215 4.170 11.375 4.790 ;
        RECT 6.895 4.170 11.375 4.330 ;
        RECT 6.895 4.170 7.055 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 8.765 4.630 9.025 4.790 ;
        RECT 4.015 4.630 5.615 4.790 ;
        RECT 5.455 4.170 5.615 4.790 ;
        RECT 5.455 4.170 6.575 4.330 ;
        RECT 6.365 4.170 6.625 4.330 ;
        RECT 6.365 4.970 6.625 5.130 ;
        RECT 6.415 4.970 8.975 5.130 ;
        RECT 8.815 4.630 8.975 5.130 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 4.975 4.170 5.135 4.790 ;
        RECT 1.615 4.170 5.135 4.330 ;
        RECT 1.615 4.170 1.775 5.130 ;
        RECT 0.175 4.970 1.775 5.130 ;
        RECT 0.175 4.630 0.335 5.130 ;
  END
END NR4D1_1
MACRO NR4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_2 0 0 ; 
  SIZE 13.260 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 4.655 5.790 ;
        RECT 3.535 5.630 4.655 5.790 ;
        RECT 3.485 5.630 3.745 5.790 ;
        RECT 4.445 5.630 4.705 5.790 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.655 0.330 3.695 0.490 ;
        RECT 0.655 0.330 0.815 3.650 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 3.695 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
    END 
  END a2
  PIN a3
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 7.805 3.490 8.065 3.650 ;
        RECT 7.855 3.490 12.335 3.650 ;
        RECT 12.125 3.490 12.385 3.650 ;
    END 
  END a3
  PIN a4
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a4
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 1.135 0.990 4.175 1.150 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 13.260 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 13.260 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 11.645 4.630 11.905 4.790 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 4.630 11.855 4.790 ;
        RECT 12.605 4.630 12.865 4.790 ;
        RECT 7.805 4.630 8.065 4.790 ;
        RECT 12.175 4.630 12.815 4.790 ;
        RECT 12.175 4.170 12.335 4.790 ;
        RECT 7.855 4.170 12.335 4.330 ;
        RECT 7.855 4.170 8.015 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 4.630 3.215 4.790 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 9.725 4.630 9.985 4.790 ;
        RECT 2.095 4.170 2.255 4.790 ;
        RECT 2.095 4.170 2.735 4.330 ;
        RECT 2.525 4.170 2.785 4.330 ;
        RECT 7.325 4.970 7.585 5.130 ;
        RECT 7.375 4.970 9.935 5.130 ;
        RECT 9.775 4.630 9.935 5.130 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 4.630 6.095 4.790 ;
  END
END NR4D1_2
#--------EOF---------

MACRO OA21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.535 0.990 4.175 1.150 ;
        RECT 3.485 0.990 3.745 1.150 ;
        RECT 0.175 0.990 0.335 4.330 ;
        RECT 0.175 4.170 1.295 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 1.135 0.330 5.135 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 4.175 5.130 ;
        RECT 4.015 4.630 4.175 5.130 ;
  END
END OA21D1
MACRO OA21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 2.575 2.530 2.735 3.170 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 2.095 2.050 3.215 2.210 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
  END
END OA21D1_1
MACRO OA21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 2.690 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 4.015 3.490 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 0.655 3.010 4.655 3.170 ;
        RECT 0.655 3.010 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 1.135 3.010 1.775 3.170 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 0.175 0.330 2.255 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END OA21D1_2
MACRO OA21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 3.485 4.630 3.745 4.790 ;
        RECT 3.055 4.630 3.695 4.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OA21D1_3
#--------EOF---------

MACRO OA21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.050 4.705 2.210 ;
        RECT 4.495 2.050 4.655 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 3.535 0.990 4.175 1.150 ;
        RECT 3.485 0.990 3.745 1.150 ;
        RECT 0.175 0.990 0.335 4.330 ;
        RECT 0.175 4.170 1.295 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 1.135 0.330 5.135 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 0.175 4.630 0.335 5.130 ;
        RECT 0.175 4.970 4.175 5.130 ;
        RECT 4.015 4.630 4.175 5.130 ;
  END
END OA21D1
MACRO OA21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_1 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.530 2.785 2.690 ;
        RECT 2.575 2.530 2.735 3.170 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 2.095 2.050 3.215 2.210 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 1.135 0.330 1.295 1.150 ;
  END
END OA21D1_1
MACRO OA21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_2 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 2.690 ;
        RECT 3.965 2.530 4.225 2.690 ;
        RECT 3.965 3.490 4.225 3.650 ;
        RECT 4.015 3.490 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.630 3.215 4.790 ;
        RECT 4.445 3.010 4.705 3.170 ;
        RECT 0.655 3.010 4.655 3.170 ;
        RECT 0.655 3.010 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 1.135 3.010 1.775 3.170 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 0.175 0.330 2.255 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END OA21D1_2
MACRO OA21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_3 0 0 ; 
  SIZE 5.440 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.630 4.225 4.790 ;
        RECT 4.015 0.990 4.175 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 5.440 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 5.440 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 3.485 4.630 3.745 4.790 ;
        RECT 3.055 4.630 3.695 4.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OA21D1_3
#--------EOF---------

MACRO OAI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1
MACRO OAI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 0.175 0.330 2.255 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END OAI21D1_1
MACRO OAI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 3.215 4.790 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.525 4.630 2.785 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1_2
MACRO OAI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 0.175 0.990 0.335 1.550 ;
        RECT 0.175 1.390 2.255 1.550 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1_3
#--------EOF---------

MACRO OAI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 2.095 0.990 2.255 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 1.135 4.170 1.295 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.070 0.335 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1
MACRO OAI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 4.630 3.215 6.050 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.175 4.630 0.335 6.050 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.055 0.070 3.215 1.150 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 0.175 0.330 2.255 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
  END
END OAI21D1_1
MACRO OAI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 0.175 0.990 0.335 4.790 ;
        RECT 0.175 4.630 3.215 4.790 ;
        RECT 2.095 0.990 2.735 1.150 ;
        RECT 2.525 0.990 2.785 1.150 ;
        RECT 2.525 4.630 2.785 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1_2
MACRO OAI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN b
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 2.690 ;
    END 
  END b
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 0.175 0.990 0.335 1.550 ;
        RECT 0.175 1.390 2.255 1.550 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.135 0.330 3.215 0.490 ;
        RECT 3.055 0.330 3.215 1.150 ;
  END
END OAI21D1_3
#--------EOF---------

MACRO OR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 0.175 3.010 2.735 3.170 ;
        RECT 0.175 3.010 0.335 4.790 ;
        RECT 1.135 0.990 1.295 3.170 ;
  END
END OR2D1
MACRO OR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.525 4.630 2.785 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END OR2D1_1
MACRO OR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 0.330 2.305 0.490 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
  END
END OR2D1_2
MACRO OR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.175 0.330 3.695 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 2.095 0.330 2.255 4.790 ;
        RECT 2.095 0.330 2.255 1.150 ;
  END
END OR2D1_3
#--------EOF---------

MACRO OR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1 0 0 ; 
  SIZE 3.740 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 3.740 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 3.740 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 0.175 3.010 2.735 3.170 ;
        RECT 0.175 3.010 0.335 4.790 ;
        RECT 1.135 0.990 1.295 3.170 ;
  END
END OR2D1
MACRO OR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_1 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.525 4.630 2.785 4.790 ;
        RECT 2.095 4.630 2.735 4.790 ;
        RECT 1.135 0.990 1.295 4.330 ;
        RECT 1.135 4.170 2.255 4.330 ;
        RECT 2.095 4.170 2.255 4.790 ;
  END
END OR2D1_1
MACRO OR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_2 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 2.045 0.330 2.305 0.490 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.990 2.255 4.790 ;
        RECT 0.175 4.630 2.255 4.790 ;
        RECT 0.175 0.990 2.255 1.150 ;
  END
END OR2D1_2
MACRO OR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_3 0 0 ; 
  SIZE 4.420 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 1.775 2.690 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.630 3.265 4.790 ;
        RECT 3.055 0.990 3.215 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 4.420 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 4.420 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 0.175 0.330 3.695 0.490 ;
        RECT 0.175 0.330 0.335 1.150 ;
        RECT 2.095 0.330 2.255 4.790 ;
        RECT 2.095 0.330 2.255 1.150 ;
  END
END OR2D1_3
#--------EOF---------

MACRO TAPCELL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL 0 0 ; 
  SIZE 2.380 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 4.700 0.600 4.860 ;
        RECT 0.390 4.700 0.550 6.050 ;
        RECT 0.820 4.700 1.080 4.860 ;
        RECT 0.870 4.700 1.030 6.050 ;
        RECT 1.300 4.700 1.560 4.860 ;
        RECT 1.350 4.700 1.510 6.050 ;
        RECT 0.000 5.970 2.380 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 0.920 0.600 1.080 ;
        RECT 0.390 0.070 0.550 1.080 ;
        RECT 0.820 0.920 1.080 1.080 ;
        RECT 0.870 0.070 1.030 1.080 ;
        RECT 1.300 0.920 1.560 1.080 ;
        RECT 1.350 0.070 1.510 1.080 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END 
  END vss 
END TAPCELL
#--------EOF---------

MACRO TAPCELL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL 0 0 ; 
  SIZE 2.380 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 4.700 0.600 4.860 ;
        RECT 0.390 4.700 0.550 6.050 ;
        RECT 0.820 4.700 1.080 4.860 ;
        RECT 0.870 4.700 1.030 6.050 ;
        RECT 1.300 4.700 1.560 4.860 ;
        RECT 1.350 4.700 1.510 6.050 ;
        RECT 0.000 5.970 2.380 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.340 0.920 0.600 1.080 ;
        RECT 0.390 0.070 0.550 1.080 ;
        RECT 0.820 0.920 1.080 1.080 ;
        RECT 0.870 0.070 1.030 1.080 ;
        RECT 1.300 0.920 1.560 1.080 ;
        RECT 1.350 0.070 1.510 1.080 ;
        RECT 0.000 -0.150 2.380 0.150 ;
    END 
  END vss 
END TAPCELL
#--------EOF---------

MACRO TIEH
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEH 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 0.655 4.630 0.815 5.130 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 0.815 1.150 ;
        RECT 0.655 0.330 0.815 1.150 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH
#--------EOF---------

MACRO TIEH
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEH 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 4.630 0.815 4.790 ;
        RECT 0.655 4.630 0.815 5.130 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 0.175 0.990 0.815 1.150 ;
        RECT 0.655 0.330 0.815 1.150 ;
        RECT 0.605 0.330 0.865 0.490 ;
  END
END TIEH
#--------EOF---------

MACRO TIEL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEL 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 0.990 0.815 1.150 ;
        RECT 0.655 0.990 0.815 1.550 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
  END
END TIEL
#--------EOF---------

MACRO TIEL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEL 0 0 ; 
  SIZE 1.700 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.175 0.990 0.815 1.150 ;
        RECT 0.655 0.990 0.815 1.550 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 4.630 1.295 6.050 ;
        RECT 0.000 5.970 1.700 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.135 0.070 1.295 1.150 ;
        RECT 0.000 -0.150 1.700 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 4.630 0.385 4.790 ;
        RECT 0.605 3.490 0.865 3.650 ;
        RECT 0.655 3.490 0.815 4.790 ;
        RECT 0.175 4.630 0.815 4.790 ;
  END
END TIEL
#--------EOF---------

MACRO XNR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 4.655 1.150 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.970 1.295 5.790 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 4.170 3.265 4.330 ;
        RECT 3.055 4.170 3.215 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 2.095 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 2.095 4.970 2.255 5.790 ;
        RECT 2.095 5.630 6.575 5.790 ;
        RECT 6.365 5.630 6.625 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.975 0.990 5.135 3.170 ;
        RECT 1.615 3.010 5.135 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 4.975 3.010 5.135 5.130 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 2.575 3.010 5.135 3.170 ;
  END
END XNR2D1
MACRO XNR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 4.970 4.175 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 0.655 0.330 3.215 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 3.055 4.970 3.215 5.790 ;
        RECT 0.655 5.630 3.215 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 3.010 3.265 3.170 ;
        RECT 3.055 3.010 3.215 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 2.095 2.530 3.215 2.690 ;
        RECT 3.055 2.530 3.215 3.170 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.975 0.990 5.135 1.550 ;
        RECT 2.575 1.390 5.135 1.550 ;
        RECT 2.575 1.390 2.735 2.210 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 4.975 1.390 5.135 5.130 ;
  END
END XNR2D1_1
MACRO XNR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 1.615 3.010 3.215 3.170 ;
        RECT 3.005 3.010 3.265 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 3.215 2.210 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 5.615 0.490 ;
        RECT 5.405 0.330 5.665 0.490 ;
        RECT 5.455 0.330 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 2.095 4.630 4.175 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 3.965 4.170 4.225 4.330 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.975 4.970 5.135 5.790 ;
        RECT 0.175 5.630 5.135 5.790 ;
        RECT 0.175 4.970 0.335 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.485 2.530 3.745 2.690 ;
        RECT 1.135 2.530 3.695 2.690 ;
        RECT 1.135 2.530 1.295 5.130 ;
        RECT 1.135 0.990 1.295 2.690 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 0.990 4.175 1.550 ;
        RECT 1.615 1.390 4.175 1.550 ;
        RECT 1.615 0.330 1.775 1.550 ;
        RECT 0.655 0.330 1.775 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 2.095 1.390 2.255 2.210 ;
        RECT 2.045 2.050 2.305 2.210 ;
        RECT 4.015 1.390 4.655 1.550 ;
        RECT 4.495 1.390 4.655 5.130 ;
        RECT 4.015 4.970 4.655 5.130 ;
  END
END XNR2D1_2
MACRO XNR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 1.615 0.330 3.695 0.490 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 3.485 4.170 3.745 4.330 ;
        RECT 0.655 4.170 3.695 4.330 ;
        RECT 0.605 4.170 0.865 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 4.655 1.150 ;
        RECT 4.495 0.330 4.655 1.150 ;
        RECT 4.495 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 4.015 0.990 4.175 4.790 ;
        RECT 2.095 4.630 4.175 4.790 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 5.455 0.990 7.055 1.150 ;
        RECT 5.455 0.990 5.615 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 4.445 4.970 4.705 5.130 ;
        RECT 0.175 4.970 4.655 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.495 4.970 7.055 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
  END
END XNR2D1_3
#--------EOF---------

MACRO XNR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 0.330 4.705 0.490 ;
        RECT 4.495 0.330 4.655 1.150 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.970 1.295 5.790 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.990 3.215 2.210 ;
        RECT 3.005 2.050 3.265 2.210 ;
        RECT 3.005 4.170 3.265 4.330 ;
        RECT 3.055 4.170 3.215 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 2.095 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 2.095 4.970 2.255 5.790 ;
        RECT 2.095 5.630 6.575 5.790 ;
        RECT 6.365 5.630 6.625 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.975 0.990 5.135 3.170 ;
        RECT 1.615 3.010 5.135 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 4.975 3.010 5.135 5.130 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 2.575 3.010 5.135 3.170 ;
  END
END XNR2D1
MACRO XNR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.495 2.530 4.655 4.330 ;
        RECT 4.445 4.170 4.705 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 2.050 3.745 2.210 ;
        RECT 3.535 2.050 3.695 3.650 ;
        RECT 3.485 3.490 3.745 3.650 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 4.970 4.175 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 4.015 0.070 4.175 1.150 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.330 3.215 1.150 ;
        RECT 0.655 0.330 3.215 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 3.055 4.970 3.215 5.790 ;
        RECT 0.655 5.630 3.215 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 3.005 3.010 3.265 3.170 ;
        RECT 3.055 3.010 3.215 4.790 ;
        RECT 2.095 4.630 3.215 4.790 ;
        RECT 2.095 4.630 2.255 5.130 ;
        RECT 2.095 0.990 2.255 2.690 ;
        RECT 2.095 2.530 3.215 2.690 ;
        RECT 3.055 2.530 3.215 3.170 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 4.975 0.990 5.135 1.550 ;
        RECT 2.575 1.390 5.135 1.550 ;
        RECT 2.575 1.390 2.735 2.210 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 4.975 1.390 5.135 5.130 ;
  END
END XNR2D1_1
MACRO XNR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 1.615 3.010 3.215 3.170 ;
        RECT 3.005 3.010 3.265 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 3.215 2.210 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 4.970 6.145 5.130 ;
        RECT 5.935 4.970 6.095 6.050 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 5.615 0.490 ;
        RECT 5.405 0.330 5.665 0.490 ;
        RECT 5.455 0.330 5.615 4.330 ;
        RECT 5.405 4.170 5.665 4.330 ;
        RECT 2.095 4.630 4.175 4.790 ;
        RECT 4.015 4.170 4.175 4.790 ;
        RECT 3.965 4.170 4.225 4.330 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.975 4.970 5.135 5.790 ;
        RECT 0.175 5.630 5.135 5.790 ;
        RECT 0.175 4.970 0.335 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 3.485 2.530 3.745 2.690 ;
        RECT 1.135 2.530 3.695 2.690 ;
        RECT 1.135 2.530 1.295 5.130 ;
        RECT 1.135 0.990 1.295 2.690 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 4.015 0.990 4.175 1.550 ;
        RECT 1.615 1.390 4.175 1.550 ;
        RECT 1.615 0.330 1.775 1.550 ;
        RECT 0.655 0.330 1.775 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 2.095 1.390 2.255 2.210 ;
        RECT 2.045 2.050 2.305 2.210 ;
        RECT 4.015 1.390 4.655 1.550 ;
        RECT 4.495 1.390 4.655 5.130 ;
        RECT 4.015 4.970 4.655 5.130 ;
  END
END XNR2D1_2
MACRO XNR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 0.330 3.745 0.490 ;
        RECT 1.615 0.330 3.695 0.490 ;
        RECT 1.565 0.330 1.825 0.490 ;
        RECT 3.485 4.170 3.745 4.330 ;
        RECT 0.655 4.170 3.695 4.330 ;
        RECT 0.605 4.170 0.865 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN zn
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END zn
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.630 2.305 4.790 ;
        RECT 2.095 0.990 4.655 1.150 ;
        RECT 4.495 0.330 4.655 1.150 ;
        RECT 4.495 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 4.015 0.990 4.175 4.790 ;
        RECT 2.095 4.630 4.175 4.790 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 5.455 0.990 7.055 1.150 ;
        RECT 5.455 0.990 5.615 3.650 ;
        RECT 5.405 3.490 5.665 3.650 ;
        RECT 4.445 4.970 4.705 5.130 ;
        RECT 0.175 4.970 4.655 5.130 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.495 4.970 7.055 5.130 ;
        RECT 0.175 4.970 0.815 5.130 ;
  END
END XNR2D1_3
#--------EOF---------

MACRO XOR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.445 4.170 4.705 4.330 ;
        RECT 2.575 4.170 4.655 4.330 ;
        RECT 2.525 4.170 2.785 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 3.535 3.490 4.175 3.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 2.210 ;
        RECT 2.095 2.050 5.135 2.210 ;
        RECT 4.925 2.050 5.185 2.210 ;
        RECT 2.095 3.490 2.255 5.130 ;
        RECT 2.045 3.490 2.305 3.650 ;
        RECT 2.045 2.050 2.305 2.210 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 2.575 0.990 3.215 1.150 ;
        RECT 2.575 0.330 2.735 1.150 ;
        RECT 0.655 0.330 2.735 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 3.055 4.970 3.215 5.790 ;
        RECT 0.655 5.630 3.215 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 3.055 0.330 5.135 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 1.615 3.010 2.735 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 2.575 3.010 5.135 3.170 ;
        RECT 4.975 3.010 5.135 5.130 ;
  END
END XOR2D1
MACRO XOR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 3.695 0.490 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 3.215 2.210 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.175 0.990 5.135 1.150 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 1.550 ;
        RECT 1.135 1.390 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 1.135 1.390 1.295 5.130 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 2.045 2.530 2.305 2.690 ;
        RECT 2.095 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 5.405 2.530 5.665 2.690 ;
        RECT 5.455 0.330 5.615 2.690 ;
        RECT 4.015 0.330 5.615 0.490 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 1.615 3.490 1.775 5.790 ;
        RECT 0.655 5.630 1.775 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 4.015 2.530 4.175 5.130 ;
  END
END XOR2D1_1
MACRO XOR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 3.695 0.490 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 0.175 0.990 4.655 1.150 ;
        RECT 4.495 0.330 4.655 1.150 ;
        RECT 4.495 0.330 7.055 0.490 ;
        RECT 6.895 0.330 7.055 1.150 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 6.895 0.990 7.055 5.130 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 1.550 ;
        RECT 1.135 1.390 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 1.135 1.390 1.295 5.130 ;
  END
END XOR2D1_2
MACRO XOR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 1.775 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.990 3.695 1.150 ;
        RECT 3.535 0.990 3.695 5.130 ;
        RECT 3.055 4.970 3.695 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 2.095 4.970 2.255 5.790 ;
        RECT 2.095 5.630 6.575 5.790 ;
        RECT 6.365 5.630 6.625 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.085 0.330 1.345 0.490 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.970 1.295 5.790 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 2.735 2.210 ;
        RECT 2.575 2.050 2.735 3.170 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 4.015 0.990 5.135 1.150 ;
        RECT 4.015 0.990 4.175 3.170 ;
        RECT 3.965 3.010 4.225 3.170 ;
        RECT 4.015 3.010 4.175 4.790 ;
        RECT 4.015 4.630 5.135 4.790 ;
        RECT 4.975 4.630 5.135 5.130 ;
  END
END XOR2D1_3
#--------EOF---------

MACRO XOR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 4.445 4.170 4.705 4.330 ;
        RECT 2.575 4.170 4.655 4.330 ;
        RECT 2.525 4.170 2.785 4.330 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 3.485 3.490 3.745 3.650 ;
        RECT 3.535 3.490 4.175 3.650 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.990 2.255 2.210 ;
        RECT 2.095 2.050 5.135 2.210 ;
        RECT 4.925 2.050 5.185 2.210 ;
        RECT 2.095 3.490 2.255 5.130 ;
        RECT 2.045 3.490 2.305 3.650 ;
        RECT 2.045 2.050 2.305 2.210 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 2.575 0.990 3.215 1.150 ;
        RECT 2.575 0.330 2.735 1.150 ;
        RECT 0.655 0.330 2.735 0.490 ;
        RECT 0.605 0.330 0.865 0.490 ;
        RECT 3.055 4.970 3.215 5.790 ;
        RECT 0.655 5.630 3.215 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 3.005 0.330 3.265 0.490 ;
        RECT 3.055 0.330 5.135 0.490 ;
        RECT 4.975 0.330 5.135 1.150 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 1.615 3.010 2.735 3.170 ;
        RECT 1.565 3.010 1.825 3.170 ;
        RECT 2.575 3.010 5.135 3.170 ;
        RECT 4.975 3.010 5.135 5.130 ;
  END
END XOR2D1
MACRO XOR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_1 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 3.695 0.490 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 3.215 2.210 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 6.845 4.630 7.105 4.790 ;
        RECT 6.895 0.990 7.055 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 0.175 0.990 5.135 1.150 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 4.975 0.990 5.135 5.130 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 1.550 ;
        RECT 1.135 1.390 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 1.135 1.390 1.295 5.130 ;
        RECT 3.965 0.990 4.225 1.150 ;
        RECT 3.965 4.970 4.225 5.130 ;
        RECT 2.045 2.530 2.305 2.690 ;
        RECT 2.095 2.530 4.655 2.690 ;
        RECT 4.445 2.530 4.705 2.690 ;
        RECT 5.405 2.530 5.665 2.690 ;
        RECT 5.455 0.330 5.615 2.690 ;
        RECT 4.015 0.330 5.615 0.490 ;
        RECT 4.015 0.330 4.175 1.150 ;
        RECT 1.565 3.490 1.825 3.650 ;
        RECT 1.615 3.490 1.775 5.790 ;
        RECT 0.655 5.630 1.775 5.790 ;
        RECT 0.605 5.630 0.865 5.790 ;
        RECT 4.015 2.530 4.175 5.130 ;
  END
END XOR2D1_1
MACRO XOR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_2 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 0.330 2.785 0.490 ;
        RECT 2.575 0.330 3.695 0.490 ;
        RECT 3.485 0.330 3.745 0.490 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 2.525 2.050 2.785 2.210 ;
        RECT 2.575 2.050 2.735 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.630 5.185 4.790 ;
        RECT 4.975 0.990 5.135 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 0.125 0.990 0.385 1.150 ;
        RECT 6.845 0.990 7.105 1.150 ;
        RECT 0.125 4.970 0.385 5.130 ;
        RECT 6.845 4.970 7.105 5.130 ;
        RECT 0.175 0.990 4.655 1.150 ;
        RECT 4.495 0.330 4.655 1.150 ;
        RECT 4.495 0.330 7.055 0.490 ;
        RECT 6.895 0.330 7.055 1.150 ;
        RECT 0.175 0.990 0.335 5.130 ;
        RECT 6.895 0.990 7.055 5.130 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.135 0.990 1.295 1.550 ;
        RECT 1.135 1.390 4.655 1.550 ;
        RECT 4.445 1.390 4.705 1.550 ;
        RECT 1.135 1.390 1.295 5.130 ;
  END
END XOR2D1_2
MACRO XOR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_3 0 0 ; 
  SIZE 7.480 BY 6.120 ; 
  SYMMETRY X Y ; 
  SITE obssite ; 
  PIN a1
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 1.565 2.530 1.825 2.690 ;
        RECT 1.615 2.530 1.775 3.170 ;
    END 
  END a1
  PIN a2
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.605 2.050 0.865 2.210 ;
        RECT 0.655 2.050 0.815 2.690 ;
    END 
  END a2
  PIN z
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER Metal1 ;
        RECT 5.885 0.990 6.145 1.150 ;
        RECT 5.885 4.630 6.145 4.790 ;
        RECT 5.935 0.990 6.095 4.790 ;
    END 
  END z
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 5.970 7.480 6.270 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER Metal1 ;
        RECT 0.000 -0.150 7.480 0.150 ;
    END 
  END vss 
  OBS
      LAYER Metal1 ;
        RECT 3.005 0.990 3.265 1.150 ;
        RECT 3.005 4.970 3.265 5.130 ;
        RECT 3.055 0.990 3.695 1.150 ;
        RECT 3.535 0.990 3.695 5.130 ;
        RECT 3.055 4.970 3.695 5.130 ;
        RECT 2.045 0.990 2.305 1.150 ;
        RECT 2.045 4.970 2.305 5.130 ;
        RECT 2.095 0.330 2.255 1.150 ;
        RECT 2.095 0.330 6.575 0.490 ;
        RECT 6.365 0.330 6.625 0.490 ;
        RECT 2.095 4.970 2.255 5.790 ;
        RECT 2.095 5.630 6.575 5.790 ;
        RECT 6.365 5.630 6.625 5.790 ;
        RECT 1.085 0.990 1.345 1.150 ;
        RECT 1.085 4.970 1.345 5.130 ;
        RECT 1.085 4.630 1.345 4.790 ;
        RECT 1.135 0.330 1.295 1.150 ;
        RECT 1.085 0.330 1.345 0.490 ;
        RECT 1.135 0.990 1.295 4.790 ;
        RECT 1.135 4.970 1.295 5.790 ;
        RECT 1.085 5.630 1.345 5.790 ;
        RECT 4.925 0.990 5.185 1.150 ;
        RECT 4.925 4.970 5.185 5.130 ;
        RECT 1.565 2.050 1.825 2.210 ;
        RECT 1.615 2.050 2.735 2.210 ;
        RECT 2.575 2.050 2.735 3.170 ;
        RECT 2.525 3.010 2.785 3.170 ;
        RECT 4.015 0.990 5.135 1.150 ;
        RECT 4.015 0.990 4.175 3.170 ;
        RECT 3.965 3.010 4.225 3.170 ;
        RECT 4.015 3.010 4.175 4.790 ;
        RECT 4.015 4.630 5.135 4.790 ;
        RECT 4.975 4.630 5.135 5.130 ;
  END
END XOR2D1_3
#--------EOF---------


END LIBRARY
