(* blackbox *)
module SARADC_CELL_INVX0_ASSW(
//`ifdef WITH_BODY
    vnw, vpw, 
//`endif
    vdd, vss, i, zn);
    input i;
    output zn;
    inout 
//`ifdef WITH_BODY
        vnw, vpw, 
//`endif
        vdd, vss;
endmodule

(* blackbox *)
module SARADC_CELL_INVX16_ASCAP(
//`ifdef WITH_BODY
    vnw, vpw, 
//`endif
    vdd, vss, i, zn);
    input i;
    output zn;
    inout 
//`ifdef WITH_BODY
        vnw, vpw, 
//`endif
        vdd, vss;
endmodule

(* blackbox *)
module SARADC_FILLTIE2(vdd, vss);
    inout vdd, vss;
endmodule

(* blackbox *)
module TIEH(z, vdd, vss);
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module TIEL(zn, vdd, vss);
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module TIEL(zn, vdd, vss);
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module INVD1(i, zn, vdd, vss);
    input i;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module INVD6(i, zn, vdd, vss);
    input i;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module INVD8(i, zn, vdd, vss);
    input i;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module OAI211D4(a1, a2, b, c, zn, vdd, vss);
    input a1, a2, b, c;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module ND2D2(a1, a2, zn, vdd, vss);
    input a1, a2;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module AN2D4(a1, a2, z, vdd, vss);
    input a1, a2;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module NR3D4(a1, a2, a3, zn, vdd, vss);
    input a1, a2, a3;
    output zn;
    inout vdd, vss;
endmodule

(* blackbox *)
module BUFFD0(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module BUFFD2(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module BUFFD4(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module BUFFD8(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module BUFFD16(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule

(* blackbox *)
module DEL4(i, z, vdd, vss);
    input i;
    output z;
    inout vdd, vss;
endmodule
