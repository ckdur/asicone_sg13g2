VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sealring
  CLASS BLOCK ;
  FOREIGN sealring ;
  ORIGIN 0.000 0.000 ;
  SIZE 1414 BY 1414 ;
  SYMMETRY X Y R90 ;
END sealring
END LIBRARY

