VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SARADC_FILL1_NOPOWER
  CLASS BLOCK ;
  FOREIGN SARADC_FILL1_NOPOWER ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.340 BY 6.120 ;
  SYMMETRY X Y R90 ;
END SARADC_FILL1_NOPOWER
END LIBRARY

