.SUBCKT sealring
.ENDS
