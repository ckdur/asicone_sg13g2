*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

.SUBCKT sg13g2_Clamp_N20N0DExt iovss pad sub
*.PININFO iovss:B pad:B
MN0 pad net2 iovss sub sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
RR1 iovss net2 1.959K $SUB=sub $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_SecondaryProtectionExt core minus pad plus sub
*.PININFO core:B minus:B pad:B plus:B
RR0 pad core 586.899 $SUB=sub $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
DD0 sub core dantenna m=1 w=640n l=3.1u a=1.984p p=7.48u
XR1 minus sub / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=640n l=4.98u a=3.187p p=11.24u
.ENDS

.SUBCKT sg13g2_Clamp_P20N0DExt iovdd iovss pad sub
*.PININFO iovdd:B iovss:B pad:B
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
XR1 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

.SUBCKT sg13g2_RCClampInverterExt in iovss out supply sub
*.PININFO in:B iovss:B out:B supply:B
MN1 iovss in iovss sub sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

.SUBCKT sg13g2_RCClampResistorExt pin1 pin2 sub
*.PININFO pin1:B pin2:B
RR29 net15 net16 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR28 net20 net21 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR27 net23 net24 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR24 net17 net18 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR23 net16 net17 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR21 net25 pin2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR20 net22 net23 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR19 net19 net20 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR17 net24 net25 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR16 net21 net22 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR15 net18 net19 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR14 net5 net6 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR13 net8 net9 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR12 net11 net12 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR11 net14 net15 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR10 net2 net3 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR9 net1 net2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR8 net13 net14 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR7 net10 net11 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR6 net7 net8 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR5 net4 net5 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR4 net12 net13 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR3 net9 net10 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR2 net6 net7 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR1 net3 net4 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR0 pin1 net1 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_Clamp_N43N43D4RExt gate pad tie sub
*.PININFO gate:I pad:B tie:B
MN0<1> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 tie sub / ptap1 r=9.999 A=65.61p Perim=32.4u w=8.1u l=8.1u
DD0 sub gate dantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

.SUBCKT sg13g2_DCNDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 anode sub / ptap1 r=5.191 A=141.253p Perim=47.54u w=11.885u l=11.885u
.ENDS

.SUBCKT sg13g2_DCPDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 guard sub / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
.ENDS

.SUBCKT sg13g2_IOPadVssExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI1 iovss vss iovss sub / sg13g2_DCNDiodeExt
XI2 vss iovdd iovss sub / sg13g2_DCPDiodeExt
XR1 iovss sub / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

.SUBCKT sg13g2_IOPadVddExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI0 net2 vdd iovss sub / sg13g2_Clamp_N43N43D4RExt
XI2 vdd net1 sub / sg13g2_RCClampResistorExt
XR1 iovss sub / ptap1 r=456.33m A=1.97n Perim=177.54u w=44.385u l=44.385u
XR0 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XI1 net1 iovss net2 vdd sub  / sg13g2_RCClampInverterExt
.ENDS

.SUBCKT sg13g2_IOPadAVDD iovdd iovss pad padres vdd vss sub
*.PININFO iovdd:B iovss:B pad:B padres:B vdd:B vss:B
XI9 iovdd iovss pad sub / sg13g2_Clamp_P20N0DExt
XI3 iovss pad iovdd sub / sg13g2_DCNDiodeExt
XI2 pad iovdd iovss sub / sg13g2_DCPDiodeExt
XI6 padres iovss pad iovdd sub / sg13g2_SecondaryProtectionExt
XI8 iovss pad sub / sg13g2_Clamp_N20N0DExt
XR1 vss sub / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS
