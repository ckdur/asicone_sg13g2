# This was copied and modified from https://github.com/IHP-GmbH/IHP-Open-PDK
# Credit to the authors

########################################################################
#
# Copyright 2023 IHP PDK Authors
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#    https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
########################################################################

VERSION 5.7 ;
#NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER contactLimit INTEGER ;
  LAYER routingPitch REAL ;
  LAYER routingGrid REAL ;
END PROPERTYDEFINITIONS

LAYER OVERLAP
   TYPE  OVERLAP ;
END OVERLAP

LAYER LOCKED
    TYPE MASTERSLICE ;
END LOCKED

LAYER LOCKED1
    TYPE MASTERSLICE ;
END LOCKED1

LAYER LOCKED2
    TYPE MASTERSLICE ;
END LOCKED2

LAYER GatPoly
  TYPE MASTERSLICE ;
END GatPoly

LAYER Cont
  TYPE CUT ;
  SPACING 0.18 ;
  WIDTH 0.16 ;
  ENCLOSURE 0 0.05 ;
  PREFERENCLOSURE 0.05 0.05 ;
  RESISTANCE 22.0 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 30 ;
    ANTENNACUMDIFFAREARATIO 10000 ;
  #PROPERTY contactLimit 10000 ;
  
END Cont

LAYER Metal1
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.48 ;
  OFFSET	0.0 ;
  WIDTH		0.16 ;
  MAXWIDTH	30 ;
  AREA		0.09 ;
  MINIMUMDENSITY        35.0 ;
  MAXIMUMDENSITY        60.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.00    1.00    10.00
  WIDTH 0.00        0.18    0.18    0.18
  WIDTH 0.30        0.18    0.22    0.22
  WIDTH 10.0        0.18    0.22    0.60 ;
  MINIMUMCUT 2 WIDTH 1.4 ;
  HEIGHT 0.930 ;
  #CURRENTDEN 0 ;
  THICKNESS 0.40 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.135 ;
  CAPACITANCE  CPERSQDIST 3.49E-05 ;
  EDGECAPACITANCE  3.16E-05 ;
  DCCURRENTDENSITY AVERAGE 1 ;

END Metal1

LAYER Via1
  TYPE	CUT ;
  RESISTANCE 20 ;
  DCCURRENTDENSITY AVERAGE 0.4 ;
  SPACING	0.22 ;
  SPACING 0.29 ADJACENTCUTS 3 WITHIN 0.311 ;
  ENCLOSURE BELOW 0.010 0.05 ;
  ENCLOSURE ABOVE 0.005 0.05 ;
  PREFERENCLOSURE 0.05 0.05 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
END Via1

LAYER Metal2
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.42 ;
  OFFSET	0.0 ;
  WIDTH		0.20 ;
  MAXWIDTH	30 ;
  MINIMUMDENSITY        35.0 ;
  MAXIMUMDENSITY        60.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.00    1.00    10.00
  WIDTH 0.00        0.21    0.21    0.21
  WIDTH 0.39        0.21    0.24    0.24
  WIDTH 10.0        0.21    0.24    0.60 ;
  MINIMUMCUT 2 WIDTH 1.4 ;
  AREA      0.144 ;
  HEIGHT 1.880 ;
  #CURRENTDEN 0 ;
  THICKNESS 0.450 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  WIREEXTENSION 0.10 ;
  RESISTANCE RPERSQ 0.103 ;
  CAPACITANCE  CPERSQDIST 1.81E-05 ;
  EDGECAPACITANCE  4.47E-05 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal2

LAYER Via2
  TYPE	CUT ;
  SPACING	0.22 ;
  WIDTH 	0.19 ;
  ENCLOSURE 0.005 0.05 ;
  PREFERENCLOSURE 0.05 0.05 ;
  RESISTANCE 20 ;
  DCCURRENTDENSITY AVERAGE 0.4 ;
  SPACING 0.29 ADJACENTCUTS 3 WITHIN 0.311 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
END Via2

LAYER Metal3
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.48 ;
  OFFSET	0.0 ;
  WIDTH		0.20 ;
  MINIMUMDENSITY        35.0 ;
  MAXIMUMDENSITY        60.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.00    1.00    10.00
  WIDTH 0.00        0.21    0.21    0.21
  WIDTH 0.39        0.21    0.24    0.24
  WIDTH 10.0        0.21    0.24    0.60 ;
  MINIMUMCUT 2 WIDTH 1.4 ;
  AREA      0.144 ;
  HEIGHT 2.880 ;
  #CURRENTDEN 0 ;
  THICKNESS 0.450 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.103 ;
  CAPACITANCE  CPERSQDIST 1.20E-05 ;
  EDGECAPACITANCE  4.48E-05 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal3

LAYER Via3
  TYPE	CUT ;
  SPACING	0.22 ;
  WIDTH 	0.19 ;
  ENCLOSURE 0.005 0.05 ;
  PREFERENCLOSURE 0.05 0.05 ;
  #RESISTANCE 0.68 ;
  RESISTANCE 20 ;
  DCCURRENTDENSITY AVERAGE 0.4 ;
  SPACING 0.29 ADJACENTCUTS 3 WITHIN 0.311 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
END Via3

LAYER Metal4
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.42 ;
  OFFSET	0.0 ;
  WIDTH		0.20 ;
  MINIMUMDENSITY        35.0 ;
  MAXIMUMDENSITY        60.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.00    1.00    10.00
  WIDTH 0.00        0.21    0.21    0.21
  WIDTH 0.39        0.21    0.24    0.24
  WIDTH 10.0        0.21    0.24    0.60 ;
  MINIMUMCUT 2 WIDTH 1.4 ;
  AREA      0.144 ;
  HEIGHT 3.88 ;
  #CURRENTDEN 0 ;
  THICKNESS 0.450 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.103 ;
  CAPACITANCE  CPERSQDIST 8.94E-06 ;
  EDGECAPACITANCE  4.50E-05 ;
  DCCURRENTDENSITY AVERAGE 2 ; #mA/um
END Metal4

LAYER Via4
  TYPE	CUT ;
  SPACING	0.22 ;
  WIDTH 0.19 ;
  ENCLOSURE 0.005 0.05 ;
  PREFERENCLOSURE 0.05 0.05 ;
  RESISTANCE 20 ;
  DCCURRENTDENSITY AVERAGE 0.4 ;
  SPACING 0.29 ADJACENTCUTS 3 WITHIN 0.311 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
END Via4

LAYER Metal5
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.48 ;
  OFFSET	0.0 ;
  WIDTH		0.20 ;
  MINIMUMDENSITY        35.0 ;
  MAXIMUMDENSITY        60.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.00    1.00    10.00
  WIDTH 0.00        0.21    0.21    0.21
  WIDTH 0.39        0.21    0.24    0.24
  WIDTH 10.0        0.21    0.24    0.60 ;
  MINIMUMCUT 2 WIDTH 1.4 ;
  AREA      0.144 ;
  HEIGHT 4.88 ;
 # CURRENTDEN 0 ;
  THICKNESS 0.450 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.103 ;
  CAPACITANCE  CPERSQDIST 7.13E-06 ;
  EDGECAPACITANCE  4.37E-05 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal5

LAYER TopVia1
  TYPE	CUT ;
  SPACING	0.42 ;
  WIDTH 	0.42 ;
  ENCLOSURE BELOW 0.1 0.1 ;
  ENCLOSURE ABOVE 0.42 0.42 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
  RESISTANCE 4.0 ;
  DCCURRENTDENSITY AVERAGE 1.4 ;
END TopVia1

LAYER TopMetal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2.28 ;
  OFFSET	1.64 ;
  WIDTH		1.64 ;
  MINIMUMDENSITY        25.0 ;
  MAXIMUMDENSITY        70.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACING 1.64 ;
  HEIGHT 6.160 ;
#  CURRENTDEN 0 ;
  THICKNESS 2.0 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.021 ;
  CAPACITANCE  CPERSQDIST 5.64E-06 ;
  EDGECAPACITANCE  5.08E-05 ;
  DCCURRENTDENSITY AVERAGE 15 ;
END TopMetal1

LAYER TopVia2
  TYPE	CUT ;
  SPACING	1.06 ;
  WIDTH 	0.9 ;
  ENCLOSURE BELOW 0.5 0.5 ;
  ENCLOSURE ABOVE 0.5 0.5 ;
  RESISTANCE 2.2 ;
  DCCURRENTDENSITY AVERAGE 10 ;
  ANTENNAAREARATIO 20 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.159 20 ) ( 0.16 80 ) ( 100 50000 ) ) ;
END TopVia2

LAYER TopMetal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		4 ;
  OFFSET	2 ;
  WIDTH		2 ;
  MINIMUMDENSITY        25.0 ;
  MAXIMUMDENSITY        70.0 ;
  DENSITYCHECKSTEP 100 ;
  DENSITYCHECKWINDOW 200 200 ;
  SPACING 2 ;
  HEIGHT 11.160 ;
#  CURRENTDEN 0 ;
  THICKNESS 3.0 ;
  ANTENNACUMAREARATIO 200 ;
  ANTENNACUMDIFFAREARATIO PWL ( ( 0 200 ) ( 0.159 200 ) ( 0.16  3200 ) ( 100 2000000 ) ) ;
  RESISTANCE RPERSQ 0.0145 ;
  CAPACITANCE  CPERSQDIST 3.23E-06 ;
  EDGECAPACITANCE  4.18E-05 ;
  DCCURRENTDENSITY AVERAGE 16 ;
END TopMetal2

#######  Via 1 Definitions ##############

Via  Via1_XX_so  DEFAULT
  RESISTANCE  20.00 ;
  LAYER  Metal1 ;
  RECT  -0.145 -0.105 0.145 0.105 ;
  LAYER  Via1 ;
  RECT  -0.095 -0.095 0.095 0.095 ;
  LAYER  Metal2 ;
  RECT  -0.145 -0.100 0.145 0.100 ;
END Via1_XX_so

Via Via1_XXE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.105 0.190 0.105 ;
    LAYER Via1 ;
        RECT -0.050 -0.095 0.140 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.100 ;
END Via1_XXE_so

Via Via1_XXW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.105 0.100 0.105 ;
    LAYER Via1 ;
        RECT -0.140 -0.095 0.050 0.095 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.100 ;
END Via1_XXW_so

Via Via1_YY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER Via1 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via1_YY_so

Via Via1_YYN_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.100 0.105 0.190 ;
    LAYER Via1 ;
        RECT -0.095 -0.050 0.095 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.190 ;
END Via1_YYN_so

Via Via1_YYS_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.190 0.105 0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.140 0.095 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.100 0.100 ;
END Via1_YYS_so

Via Via1_XY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.145 -0.105 0.145 0.105 ;
    LAYER Via1 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via1_XY_so

Via Via1_XYNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.080 0.100 0.150 ;
    LAYER Via1 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.150 -0.100 0.100 0.190 ;
END Via1_XYNW_so

Via Via1_XYNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.080 0.190 0.150 ;
    LAYER Via1 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.150 0.190 ;
END Via1_XYNE_so

Via Via1_XYSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.150 0.190 0.080 ;
    LAYER Via1 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.150 0.100 ;
END Via1_XYSE_so

Via Via1_XYSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.150 0.100 0.080 ;
    LAYER Via1 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.150 -0.190 0.100 0.100 ;
END Via1_XYSW_so

Via Via1_YX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER Via1 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via1_YX_so

Via Via1_YXNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.150 -0.100 0.080 0.190 ;
    LAYER Via1 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.150 ;
END Via1_YXNW_so

Via Via1_YXNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.080 -0.100 0.150 0.190 ;
    LAYER Via1 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.150 ;
END Via1_YXNE_so

Via Via1_YXSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.080 -0.190 0.150 0.100 ;
    LAYER Via1 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.150 0.190 0.100 ;
END Via1_YXSE_so

Via Via1_YXSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.150 -0.190 0.080 0.100 ;
    LAYER Via1 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.190 -0.150 0.100 0.100 ;
END Via1_YXSW_so

##############

Via Via1_NE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.190 0.190 ;
    LAYER Via1 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.190 ;
END Via1_NE_eo

Via Via1_NW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.100 0.100 0.190 ;
    LAYER Via1 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.190 ;
END Via1_NW_eo

Via Via1_SE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.190 0.190 0.100 ;
    LAYER Via1 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.190 0.100 ;
END Via1_SE_eo

Via Via1_SW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.190 0.100 0.100 ;
    LAYER Via1 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.190 -0.190 0.100 0.100 ;
END Via1_SW_eo

##############

Via Via1_NE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.250 0.250 ;
    LAYER Via1 ;
        RECT -0.020 -0.020 0.170 0.170 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.250 0.250 ;
END Via1_NE_beo

Via Via1_NW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.250 -0.100 0.100 0.250 ;
    LAYER Via1 ;
        RECT -0.170 -0.020 0.020 0.170 ;
    LAYER Metal2 ;
        RECT -0.250 -0.100 0.100 0.250 ;
END Via1_NW_beo

Via Via1_SE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.250 0.250 0.100 ;
    LAYER Via1 ;
        RECT -0.020 -0.170 0.170 0.020 ;
    LAYER Metal2 ;
        RECT -0.100 -0.250 0.250 0.100 ;
END Via1_SE_beo

Via Via1_SW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal1 ;
        RECT -0.250 -0.250 0.100 0.100 ;
    LAYER Via1 ;
        RECT -0.170 -0.170 0.020 0.020 ;
    LAYER Metal2 ;
        RECT -0.250 -0.250 0.100 0.100 ;
END Via1_SW_beo

##############

Via Via1_DV1E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.105 0.600 0.105 ;
    LAYER Via1 ;
        RECT -0.050 -0.095 0.140 0.095 ;
        RECT  0.360 -0.095 0.550 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.600 0.100 ;
END Via1_DV1E_so

Via Via1_DV1W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.600 -0.105  0.100 0.105 ;
    LAYER Via1 ;
        RECT -0.550 -0.095 -0.360 0.095 ;
        RECT -0.140 -0.095  0.050 0.095 ;
    LAYER Metal2 ;
        RECT -0.600 -0.100  0.100 0.100 ;
END Via1_DV1W_so

Via Via1_DV1S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.600 0.105  0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.140 0.095  0.050 ;
        RECT -0.095 -0.550 0.095 -0.360 ;
    LAYER Metal2 ;
        RECT -0.100 -0.600 0.100  0.100 ;
END Via1_DV1S_so

Via Via1_DV1SM_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.560 0.105  0.140 ;
    LAYER Via1 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.560 0.100  0.140 ;
END Via1_DV1SM_so

Via Via1_DV1N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.100 0.105 0.600 ;
    LAYER Via1 ;
        RECT -0.095 -0.050 0.095 0.140 ;
        RECT -0.095  0.360 0.095 0.550 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.600 ;
END Via1_DV1N_so

Via Via1_DV1NM_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.140 0.105  0.560 ;
    LAYER Via1 ;
        RECT -0.095  0.320 0.095  0.510 ;
        RECT -0.095 -0.090 0.095  0.100 ;
    LAYER Metal2 ;
        RECT -0.100 -0.140 0.100  0.560 ;
END Via1_DV1NM_so

Via Via1_DV2E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.140 -0.105 0.560 0.105 ;
    LAYER Via1 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via1_DV2E_so

Via Via1_DV2EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.140 -0.100 0.560 0.150 ;
    LAYER Via1 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via1_DV2EN_so

Via Via1_DV2ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.140 -0.150 0.560 0.100 ;
    LAYER Via1 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via1_DV2ES_so

Via Via1_DV2W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.560 -0.105  0.140 0.105 ;
    LAYER Via1 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal2 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via1_DV2W_so

Via Via1_DV2WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.560 -0.100  0.140 0.150 ;
    LAYER Via1 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via1_DV2WN_so

Via Via1_DV2WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.560 -0.150  0.140 0.100 ;
    LAYER Via1 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal2 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via1_DV2WS_so

Via Via1_DV2S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.560 0.100  0.140 ;
END Via1_DV2S_so

Via Via1_DV2SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via1 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.560 0.150  0.140 ;
END Via1_DV2SE_so

Via Via1_DV2SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via1 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal2 ;
        RECT -0.150 -0.560 0.100  0.140 ;
END Via1_DV2SW_so

Via Via1_DV2N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via1 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.140 0.100 0.560 ;
END Via1_DV2N_so

Via Via1_DV2NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via1 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.140 0.150 0.560 ;
END Via1_DV2NE_so

Via Via1_DV2NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via1 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal2 ;
        RECT -0.150 -0.140 0.100 0.560 ;
END Via1_DV2NW_so

##############

Via Via1_DV3E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.520 0.145 ;
    LAYER Via1 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal1 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via1_DV3E_so

Via Via1_DV3EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.190 ;
    LAYER Via1 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via1_DV3EN_so

Via Via1_DV3ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.520 0.100 ;
    LAYER Via1 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal1 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via1_DV3ES_so

Via Via1_DV3W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.520 -0.145  0.100 0.145 ;
    LAYER Via1 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal1 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via1_DV3W_so

Via Via1_DV3WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.190 ;
    LAYER Via1 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal1 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via1_DV3WN_so

Via Via1_DV3WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.520 -0.190  0.100 0.100 ;
    LAYER Via1 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal1 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via1_DV3WS_so

Via Via1_DV3S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal1 ;
        RECT -0.145 -0.520 0.145  0.100 ;
END Via1_DV3S_so

Via Via1_DV3SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via1 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal1 ;
        RECT -0.100 -0.520 0.190  0.100 ;
END Via1_DV3SE_so

Via Via1_DV3SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via1 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal1 ;
        RECT -0.190 -0.520 0.100  0.100 ;
END Via1_DV3SW_so

Via Via1_DV3N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via1 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal1 ;
        RECT -0.145 -0.100 0.145 0.520 ;
END Via1_DV3N_so

Via Via1_DV3NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via1 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.190 0.520 ;
END Via1_DV3NE_so

Via Via1_DV3NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via1 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal1 ;
        RECT -0.190 -0.100 0.100 0.520 ;
END Via1_DV3NW_so

##############

Via Via1_DV1E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.105 0.660 0.105 ;
    LAYER Via1 ;
        RECT -0.020 -0.095 0.170 0.095 ;
        RECT  0.390 -0.095 0.580 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.660 0.100 ;
END Via1_DV1E_eo

Via Via1_DV1W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.660 -0.105  0.100 0.105 ;
    LAYER Via1 ;
        RECT -0.580 -0.095 -0.390 0.095 ;
        RECT -0.170 -0.095  0.020 0.095 ;
    LAYER Metal2 ;
        RECT -0.660 -0.100  0.100 0.100 ;
END Via1_DV1W_eo

Via Via1_DV1S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.660 0.105  0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.170 0.095  0.020 ;
        RECT -0.095 -0.580 0.095 -0.390 ;
    LAYER Metal2 ;
        RECT -0.100 -0.660 0.100  0.100 ;
END Via1_DV1S_eo

Via Via1_DV1N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.105 -0.100 0.105 0.660 ;
    LAYER Via1 ;
        RECT -0.095 -0.020 0.095 0.170 ;
        RECT -0.095  0.390 0.095 0.580 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.660 ;
END Via1_DV1N_eo

Via Via1_DV2E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.170 -0.105 0.590 0.105 ;
    LAYER Via1 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.175 0.520 0.175 ;
END Via1_DV2E_eo

Via Via1_DV2EN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.170 -0.100 0.590 0.180 ;
    LAYER Via1 ;
        RECT -0.090 -0.020 0.100 0.170 ;
        RECT  0.320 -0.020 0.510 0.170 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.250 ;
END Via1_DV2EN_eo

Via Via1_DV2ES_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.170 -0.180 0.590 0.100 ;
    LAYER Via1 ;
        RECT -0.090 -0.170 0.100 0.020 ;
        RECT  0.320 -0.170 0.510 0.020 ;
    LAYER Metal2 ;
        RECT -0.100 -0.250 0.520 0.100 ;
END Via1_DV2ES_eo

Via Via1_DV2W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.590 -0.105  0.170 0.105 ;
    LAYER Via1 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal2 ;
        RECT -0.520 -0.175  0.100 0.175 ;
END Via1_DV2W_eo

Via Via1_DV2WN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.590 -0.100  0.170 0.180 ;
    LAYER Via1 ;
        RECT -0.510 -0.020 -0.320 0.170 ;
        RECT -0.100 -0.020  0.090 0.170 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.250 ;
END Via1_DV2WN_eo

Via Via1_DV2WS_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.590 -0.180  0.170 0.100 ;
    LAYER Via1 ;
        RECT -0.510 -0.170 -0.320 0.020 ;
        RECT -0.100 -0.170  0.090 0.020 ;
    LAYER Metal2 ;
        RECT -0.520 -0.250  0.100 0.100 ;
END Via1_DV2WS_eo

Via Via1_DV2S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.175 -0.520 0.175  0.100 ;
    LAYER Via1 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.590 0.100  0.170 ;
END Via1_DV2S_eo

Via Via1_DV2SE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.520 0.250  0.100 ;
    LAYER Via1 ;
        RECT -0.020 -0.100 0.170  0.090 ;
        RECT -0.020 -0.510 0.170 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.590 0.220  0.170 ;
END Via1_DV2SE_eo

Via Via1_DV2SW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.250 -0.520 0.100  0.100 ;
    LAYER Via1 ;
        RECT -0.170 -0.100 0.020  0.090 ;
        RECT -0.170 -0.510 0.020 -0.320 ;
    LAYER Metal2 ;
        RECT -0.220 -0.590 0.100  0.170 ;
END Via1_DV2SW_eo

Via Via1_DV2N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.175 -0.100 0.175 0.520 ;
    LAYER Via1 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.170 0.100 0.590 ;
END Via1_DV2N_eo

Via Via1_DV2NE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.250 0.520 ;
    LAYER Via1 ;
        RECT -0.020 -0.090 0.170 0.100 ;
        RECT -0.020  0.320 0.170 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.170 0.220 0.590 ;
END Via1_DV2NE_eo

Via Via1_DV2NW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.250 -0.100 0.100 0.520 ;
    LAYER Via1 ;
        RECT -0.170 -0.090 0.020 0.100 ;
        RECT -0.170  0.320 0.020 0.510 ;
    LAYER Metal2 ;
        RECT -0.220 -0.170 0.100 0.590 ;
END Via1_DV2NW_eo

##############

Via Via1_DV1EN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.100 0.660 0.190 ;
    LAYER Via1 ;
        RECT -0.020 -0.050 0.170 0.140 ;
        RECT  0.390 -0.050 0.580 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.660 0.190 ;
END Via1_DV1EN_beo

Via Via1_DV1ES_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.190 0.660 0.100 ;
    LAYER Via1 ;
        RECT -0.020 -0.140 0.170 0.050 ;
        RECT  0.390 -0.140 0.580 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.660 0.100 ;
END Via1_DV1ES_beo

Via Via1_DV1WN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.660 -0.100  0.100 0.190 ;
    LAYER Via1 ;
        RECT -0.580 -0.050 -0.390 0.140 ;
        RECT -0.170 -0.050  0.020 0.140 ;
    LAYER Metal2 ;
        RECT -0.660 -0.100  0.100 0.190 ;
END Via1_DV1WN_beo

Via Via1_DV1WS_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.660 -0.190  0.100 0.100 ;
    LAYER Via1 ;
        RECT -0.580 -0.140 -0.390 0.050 ;
        RECT -0.170 -0.140  0.020 0.050 ;
    LAYER Metal2 ;
        RECT -0.660 -0.190  0.100 0.100 ;
END Via1_DV1WS_beo

Via Via1_DV1SE_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.100 -0.660 0.190  0.100 ;
    LAYER Via1 ;
        RECT -0.050 -0.170 0.140  0.020 ;
        RECT -0.050 -0.580 0.140 -0.390 ;
    LAYER Metal2 ;
        RECT -0.100 -0.660 0.190  0.100 ;
END Via1_DV1SE_beo

Via Via1_DV1SW_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal1 ;
        RECT -0.190 -0.660 0.100  0.100 ;
    LAYER Via1 ;
        RECT -0.140 -0.170 0.050  0.020 ;
        RECT -0.140 -0.580 0.050 -0.390 ;
    LAYER Metal2 ;
        RECT -0.190 -0.660 0.100  0.100 ;
END Via1_DV1SW_beo

######### Via 2 Definitions ##############
Via Via2_XX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via2_XX_so

Via Via2_XXE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.095 0.140 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.100 ;
END Via2_XXE_so

Via Via2_XXW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.095 0.050 0.095 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.100 ;
END Via2_XXW_so

Via Via2_YY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via2 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via2_YY_so

Via Via2_YYN_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.190 ;
    LAYER Via2 ;
        RECT -0.095 -0.050 0.095 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.190 ;
END Via2_YYN_so

Via Via2_YYS_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.140 0.095 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.100 0.100 ;
END Via2_YYS_so

Via Via2_XY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via2_XY_so

Via Via2_XYNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.150 ;
    LAYER Via2 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.150 -0.100 0.100 0.190 ;
END Via2_XYNW_so

Via Via2_XYNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.150 ;
    LAYER Via2 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.150 0.190 ;
END Via2_XYNE_so

Via Via2_XYSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.150 0.190 0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.150 0.100 ;
END Via2_XYSE_so

Via Via2_XYSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.150 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.150 -0.190 0.100 0.100 ;
END Via2_XYSW_so

Via Via2_YX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via2 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal2 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via2_YX_so

Via Via2_YXNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.150 -0.100 0.100 0.190 ;
    LAYER Via2 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.150 ;
END Via2_YXNW_so

Via Via2_YXNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.150 0.190 ;
    LAYER Via2 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.150 ;
END Via2_YXNE_so

Via Via2_YXSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.150 0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.150 0.190 0.100 ;
END Via2_YXSE_so

Via Via2_YXSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.150 -0.190 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.190 -0.150 0.100 0.100 ;
END Via2_YXSW_so

##############

Via Via2_NE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.190 ;
    LAYER Via2 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.190 ;
END Via2_NE_eo

Via Via2_NW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.190 ;
    LAYER Via2 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.190 ;
END Via2_NW_eo

Via Via2_SE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.190 0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.190 0.100 ;
END Via2_SE_eo

Via Via2_SW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.190 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal2 ;
        RECT -0.190 -0.190 0.100 0.100 ;
END Via2_SW_eo

##############

Via Via2_NE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.250 0.250 ;
    LAYER Via2 ;
        RECT -0.020 -0.020 0.170 0.170 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.250 0.250 ;
END Via2_NE_beo

Via Via2_NW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.100 0.100 0.250 ;
    LAYER Via2 ;
        RECT -0.170 -0.020 0.020 0.170 ;
    LAYER Metal2 ;
        RECT -0.250 -0.100 0.100 0.250 ;
END Via2_NW_beo

Via Via2_SE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.250 0.250 0.100 ;
    LAYER Via2 ;
        RECT -0.020 -0.170 0.170 0.020 ;
    LAYER Metal2 ;
        RECT -0.100 -0.250 0.250 0.100 ;
END Via2_SE_beo

Via Via2_SW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.250 0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.170 -0.170 0.020 0.020 ;
    LAYER Metal2 ;
        RECT -0.250 -0.250 0.100 0.100 ;
END Via2_SW_beo

##############

Via Via2_DV1E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.600 0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.095 0.140 0.095 ;
        RECT  0.360 -0.095 0.550 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.600 0.100 ;
END Via2_DV1E_so

Via Via2_DV1W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.600 -0.100  0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.550 -0.095 -0.360 0.095 ;
        RECT -0.140 -0.095  0.050 0.095 ;
    LAYER Metal2 ;
        RECT -0.600 -0.100  0.100 0.100 ;
END Via2_DV1W_so

Via Via2_DV1S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.600 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.140 0.095  0.050 ;
        RECT -0.095 -0.550 0.095 -0.360 ;
    LAYER Metal2 ;
        RECT -0.100 -0.600 0.100  0.100 ;
END Via2_DV1S_so

Via Via2_DV1N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.600 ;
    LAYER Via2 ;
        RECT -0.095 -0.050 0.095 0.140 ;
        RECT -0.095  0.360 0.095 0.550 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.600 ;
END Via2_DV1N_so

Via Via2_DV2E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.100 0.560 0.100 ;
    LAYER Via2 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via2_DV2E_so

Via Via2_DV2EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.100 0.560 0.150 ;
    LAYER Via2 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via2_DV2EN_so

Via Via2_DV2ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.150 0.560 0.100 ;
    LAYER Via2 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via2_DV2ES_so

Via Via2_DV2W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.100  0.140 0.100 ;
    LAYER Via2 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal2 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via2_DV2W_so

Via Via2_DV2WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.100  0.140 0.150 ;
    LAYER Via2 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via2_DV2WN_so

Via Via2_DV2WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.150  0.140 0.100 ;
    LAYER Via2 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal2 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via2_DV2WS_so

Via Via2_DV2S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.560 0.100  0.140 ;
END Via2_DV2S_so

Via Via2_DV2SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.560 0.150  0.140 ;
END Via2_DV2SE_so

Via Via2_DV2SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal2 ;
        RECT -0.150 -0.560 0.100  0.140 ;
END Via2_DV2SW_so

Via Via2_DV2N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via2 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.140 0.100 0.560 ;
END Via2_DV2N_so

Via Via2_DV2NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via2 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.140 0.150 0.560 ;
END Via2_DV2NE_so

Via Via2_DV2NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via2 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal2 ;
        RECT -0.150 -0.140 0.100 0.560 ;
END Via2_DV2NW_so

##############

Via Via2_DV3E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.520 0.145 ;
    LAYER Via2 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via2_DV3E_so

Via Via2_DV3EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.520 0.190 ;
    LAYER Via2 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via2_DV3EN_so

Via Via2_DV3ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.520 0.100 ;
    LAYER Via2 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via2_DV3ES_so

Via Via2_DV3W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.520 -0.145  0.100 0.145 ;
    LAYER Via2 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal2 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via2_DV3W_so

Via Via2_DV3WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.520 -0.100  0.100 0.190 ;
    LAYER Via2 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via2_DV3WN_so

Via Via2_DV3WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.520 -0.190  0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal2 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via2_DV3WS_so

Via Via2_DV3S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.145 -0.520 0.145  0.100 ;
END Via2_DV3S_so

Via Via2_DV3SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.520 0.190  0.100 ;
END Via2_DV3SE_so

Via Via2_DV3SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal2 ;
        RECT -0.190 -0.520 0.100  0.100 ;
END Via2_DV3SW_so

Via Via2_DV3N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via2 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal2 ;
        RECT -0.145 -0.100 0.145 0.520 ;
END Via2_DV3N_so

Via Via2_DV3NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via2 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.190 0.520 ;
END Via2_DV3NE_so

Via Via2_DV3NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via2 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal2 ;
        RECT -0.190 -0.100 0.100 0.520 ;
END Via2_DV3NW_so

##############

Via Via2_DV1E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.660 0.100 ;
    LAYER Via2 ;
        RECT -0.020 -0.095 0.170 0.095 ;
        RECT  0.390 -0.095 0.580 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.660 0.100 ;
END Via2_DV1E_eo

Via Via2_DV1W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.100  0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.580 -0.095 -0.390 0.095 ;
        RECT -0.170 -0.095  0.020 0.095 ;
    LAYER Metal2 ;
        RECT -0.660 -0.100  0.100 0.100 ;
END Via2_DV1W_eo

Via Via2_DV1S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.660 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.170 0.095  0.020 ;
        RECT -0.095 -0.580 0.095 -0.390 ;
    LAYER Metal2 ;
        RECT -0.100 -0.660 0.100  0.100 ;
END Via2_DV1S_eo

Via Via2_DV1N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.660 ;
    LAYER Via2 ;
        RECT -0.095 -0.020 0.095 0.170 ;
        RECT -0.095  0.390 0.095 0.580 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.100 0.660 ;
END Via2_DV1N_eo

Via Via2_DV2E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.100 0.590 0.100 ;
    LAYER Via2 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal2 ;
        RECT -0.100 -0.175 0.520 0.175 ;
END Via2_DV2E_eo

Via Via2_DV2EN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.100 0.590 0.180 ;
    LAYER Via2 ;
        RECT -0.090 -0.020 0.100 0.170 ;
        RECT  0.320 -0.020 0.510 0.170 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.520 0.250 ;
END Via2_DV2EN_eo

Via Via2_DV2ES_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.180 0.590 0.100 ;
    LAYER Via2 ;
        RECT -0.090 -0.170 0.100 0.020 ;
        RECT  0.320 -0.170 0.510 0.020 ;
    LAYER Metal2 ;
        RECT -0.100 -0.250 0.520 0.100 ;
END Via2_DV2ES_eo

Via Via2_DV2W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.100  0.170 0.100 ;
    LAYER Via2 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal2 ;
        RECT -0.520 -0.175  0.100 0.175 ;
END Via2_DV2W_eo

Via Via2_DV2WN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.100  0.170 0.180 ;
    LAYER Via2 ;
        RECT -0.510 -0.020 -0.320 0.170 ;
        RECT -0.100 -0.020  0.090 0.170 ;
    LAYER Metal2 ;
        RECT -0.520 -0.100  0.100 0.250 ;
END Via2_DV2WN_eo

Via Via2_DV2WS_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.180  0.170 0.100 ;
    LAYER Via2 ;
        RECT -0.510 -0.170 -0.320 0.020 ;
        RECT -0.100 -0.170  0.090 0.020 ;
    LAYER Metal2 ;
        RECT -0.520 -0.250  0.100 0.100 ;
END Via2_DV2WS_eo

Via Via2_DV2S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.175 -0.520 0.175  0.100 ;
    LAYER Via2 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.590 0.100  0.170 ;
END Via2_DV2S_eo

Via Via2_DV2SE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.250  0.100 ;
    LAYER Via2 ;
        RECT -0.020 -0.100 0.170  0.090 ;
        RECT -0.020 -0.510 0.170 -0.320 ;
    LAYER Metal2 ;
        RECT -0.100 -0.590 0.220  0.170 ;
END Via2_DV2SE_eo

Via Via2_DV2SW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.520 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.170 -0.100 0.020  0.090 ;
        RECT -0.170 -0.510 0.020 -0.320 ;
    LAYER Metal2 ;
        RECT -0.220 -0.590 0.100  0.170 ;
END Via2_DV2SW_eo

Via Via2_DV2N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.175 -0.100 0.175 0.520 ;
    LAYER Via2 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.170 0.100 0.590 ;
END Via2_DV2N_eo

Via Via2_DV2NE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.250 0.520 ;
    LAYER Via2 ;
        RECT -0.020 -0.090 0.170 0.100 ;
        RECT -0.020  0.320 0.170 0.510 ;
    LAYER Metal2 ;
        RECT -0.100 -0.170 0.220 0.590 ;
END Via2_DV2NE_eo

Via Via2_DV2NW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.100 0.100 0.520 ;
    LAYER Via2 ;
        RECT -0.170 -0.090 0.020 0.100 ;
        RECT -0.170  0.320 0.020 0.510 ;
    LAYER Metal2 ;
        RECT -0.220 -0.170 0.100 0.590 ;
END Via2_DV2NW_eo

##############

Via Via2_DV1EN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.660 0.190 ;
    LAYER Via2 ;
        RECT -0.020 -0.050 0.170 0.140 ;
        RECT  0.390 -0.050 0.580 0.140 ;
    LAYER Metal2 ;
        RECT -0.100 -0.100 0.660 0.190 ;
END Via2_DV1EN_beo

Via Via2_DV1ES_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.660 0.100 ;
    LAYER Via2 ;
        RECT -0.020 -0.140 0.170 0.050 ;
        RECT  0.390 -0.140 0.580 0.050 ;
    LAYER Metal2 ;
        RECT -0.100 -0.190 0.660 0.100 ;
END Via2_DV1ES_beo

Via Via2_DV1WN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.100  0.100 0.190 ;
    LAYER Via2 ;
        RECT -0.580 -0.050 -0.390 0.140 ;
        RECT -0.170 -0.050  0.020 0.140 ;
    LAYER Metal2 ;
        RECT -0.660 -0.100  0.100 0.190 ;
END Via2_DV1WN_beo

Via Via2_DV1WS_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.190  0.100 0.100 ;
    LAYER Via2 ;
        RECT -0.580 -0.140 -0.390 0.050 ;
        RECT -0.170 -0.140  0.020 0.050 ;
    LAYER Metal2 ;
        RECT -0.660 -0.190  0.100 0.100 ;
END Via2_DV1WS_beo

Via Via2_DV1SE_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.660 0.190  0.100 ;
    LAYER Via2 ;
        RECT -0.050 -0.170 0.140  0.020 ;
        RECT -0.050 -0.580 0.140 -0.390 ;
    LAYER Metal2 ;
        RECT -0.100 -0.660 0.190  0.100 ;
END Via2_DV1SE_beo

Via Via2_DV1SW_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.660 0.100  0.100 ;
    LAYER Via2 ;
        RECT -0.140 -0.170 0.050  0.020 ;
        RECT -0.140 -0.580 0.050 -0.390 ;
    LAYER Metal2 ;
        RECT -0.190 -0.660 0.100  0.100 ;
END Via2_DV1SW_beo

######### Via 3 Definitions ######################
Via Via3_XX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via3_XX_so

Via Via3_XXE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.095 0.140 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.100 ;
END Via3_XXE_so

Via Via3_XXW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.095 0.050 0.095 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.100 ;
END Via3_XXW_so

Via Via3_YY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via3 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via3_YY_so

Via Via3_YYN_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.190 ;
    LAYER Via3 ;
        RECT -0.095 -0.050 0.095 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.190 ;
END Via3_YYN_so

Via Via3_YYS_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.140 0.095 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.100 0.100 ;
END Via3_YYS_so

Via Via3_XY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via3_XY_so

Via Via3_XYNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.150 ;
    LAYER Via3 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.150 -0.100 0.100 0.190 ;
END Via3_XYNW_so

Via Via3_XYNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.150 ;
    LAYER Via3 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.150 0.190 ;
END Via3_XYNE_so

Via Via3_XYSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.150 0.190 0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.150 0.100 ;
END Via3_XYSE_so

Via Via3_XYSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.150 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.150 -0.190 0.100 0.100 ;
END Via3_XYSW_so

Via Via3_YX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via3 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via3_YX_so

Via Via3_YXNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.150 -0.100 0.100 0.190 ;
    LAYER Via3 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.150 ;
END Via3_YXNW_so

Via Via3_YXNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.150 0.190 ;
    LAYER Via3 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.150 ;
END Via3_YXNE_so

Via Via3_YXSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.150 0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.150 0.190 0.100 ;
END Via3_YXSE_so

Via Via3_YXSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.150 -0.190 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.190 -0.150 0.100 0.100 ;
END Via3_YXSW_so

##############

Via Via3_NE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.190 ;
    LAYER Via3 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.190 ;
END Via3_NE_eo

Via Via3_NW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.190 ;
    LAYER Via3 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.190 ;
END Via3_NW_eo

Via Via3_SE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.190 0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.190 0.100 ;
END Via3_SE_eo

Via Via3_SW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.190 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.190 -0.190 0.100 0.100 ;
END Via3_SW_eo

##############

Via Via3_NE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.250 0.250 ;
    LAYER Via3 ;
        RECT -0.020 -0.020 0.170 0.170 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.250 0.250 ;
END Via3_NE_beo

Via Via3_NW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.100 0.100 0.250 ;
    LAYER Via3 ;
        RECT -0.170 -0.020 0.020 0.170 ;
    LAYER Metal4 ;
        RECT -0.250 -0.100 0.100 0.250 ;
END Via3_NW_beo

Via Via3_SE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.250 0.250 0.100 ;
    LAYER Via3 ;
        RECT -0.020 -0.170 0.170 0.020 ;
    LAYER Metal4 ;
        RECT -0.100 -0.250 0.250 0.100 ;
END Via3_SE_beo

Via Via3_SW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.250 0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.170 -0.170 0.020 0.020 ;
    LAYER Metal4 ;
        RECT -0.250 -0.250 0.100 0.100 ;
END Via3_SW_beo

##############

Via Via3_DV1E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.600 0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.095 0.140 0.095 ;
        RECT  0.360 -0.095 0.550 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.600 0.100 ;
END Via3_DV1E_so

Via Via3_DV1W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.600 -0.100  0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.550 -0.095 -0.360 0.095 ;
        RECT -0.140 -0.095  0.050 0.095 ;
    LAYER Metal4 ;
        RECT -0.600 -0.100  0.100 0.100 ;
END Via3_DV1W_so

Via Via3_DV1S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.600 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.140 0.095  0.050 ;
        RECT -0.095 -0.550 0.095 -0.360 ;
    LAYER Metal4 ;
        RECT -0.100 -0.600 0.100  0.100 ;
END Via3_DV1S_so

Via Via3_DV1N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.600 ;
    LAYER Via3 ;
        RECT -0.095 -0.050 0.095 0.140 ;
        RECT -0.095  0.360 0.095 0.550 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.600 ;
END Via3_DV1N_so

Via Via3_DV2E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.100 0.560 0.100 ;
    LAYER Via3 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via3_DV2E_so

Via Via3_DV2EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.100 0.560 0.150 ;
    LAYER Via3 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via3_DV2EN_so

Via Via3_DV2ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.140 -0.150 0.560 0.100 ;
    LAYER Via3 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via3_DV2ES_so

Via Via3_DV2W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.100  0.140 0.100 ;
    LAYER Via3 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal4 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via3_DV2W_so

Via Via3_DV2WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.100  0.140 0.150 ;
    LAYER Via3 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via3_DV2WN_so

Via Via3_DV2WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.560 -0.150  0.140 0.100 ;
    LAYER Via3 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal4 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via3_DV2WS_so

Via Via3_DV2S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.560 0.100  0.140 ;
END Via3_DV2S_so

Via Via3_DV2SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.560 0.150  0.140 ;
END Via3_DV2SE_so

Via Via3_DV2SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal4 ;
        RECT -0.150 -0.560 0.100  0.140 ;
END Via3_DV2SW_so

Via Via3_DV2N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via3 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.140 0.100 0.560 ;
END Via3_DV2N_so

Via Via3_DV2NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via3 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.140 0.150 0.560 ;
END Via3_DV2NE_so

Via Via3_DV2NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via3 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal4 ;
        RECT -0.150 -0.140 0.100 0.560 ;
END Via3_DV2NW_so

##############

Via Via3_DV3E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.520 0.145 ;
    LAYER Via3 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal3 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via3_DV3E_so

Via Via3_DV3EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.190 ;
    LAYER Via3 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via3_DV3EN_so

Via Via3_DV3ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.520 0.100 ;
    LAYER Via3 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via3_DV3ES_so

Via Via3_DV3W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.520 -0.145  0.100 0.145 ;
    LAYER Via3 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal3 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via3_DV3W_so

Via Via3_DV3WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.190 ;
    LAYER Via3 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal3 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via3_DV3WN_so

Via Via3_DV3WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.520 -0.190  0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal3 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via3_DV3WS_so

Via Via3_DV3S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal3 ;
        RECT -0.145 -0.520 0.145  0.100 ;
END Via3_DV3S_so

Via Via3_DV3SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.190  0.100 ;
END Via3_DV3SE_so

Via Via3_DV3SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal3 ;
        RECT -0.190 -0.520 0.100  0.100 ;
END Via3_DV3SW_so

Via Via3_DV3N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via3 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal3 ;
        RECT -0.145 -0.100 0.145 0.520 ;
END Via3_DV3N_so

Via Via3_DV3NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via3 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.190 0.520 ;
END Via3_DV3NE_so

Via Via3_DV3NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via3 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal3 ;
        RECT -0.190 -0.100 0.100 0.520 ;
END Via3_DV3NW_so

##############

Via Via3_DV1E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.660 0.100 ;
    LAYER Via3 ;
        RECT -0.020 -0.095 0.170 0.095 ;
        RECT  0.390 -0.095 0.580 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.660 0.100 ;
END Via3_DV1E_eo

Via Via3_DV1W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.100  0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.580 -0.095 -0.390 0.095 ;
        RECT -0.170 -0.095  0.020 0.095 ;
    LAYER Metal4 ;
        RECT -0.660 -0.100  0.100 0.100 ;
END Via3_DV1W_eo

Via Via3_DV1S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.660 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.170 0.095  0.020 ;
        RECT -0.095 -0.580 0.095 -0.390 ;
    LAYER Metal4 ;
        RECT -0.100 -0.660 0.100  0.100 ;
END Via3_DV1S_eo

Via Via3_DV1N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.100 0.660 ;
    LAYER Via3 ;
        RECT -0.095 -0.020 0.095 0.170 ;
        RECT -0.095  0.390 0.095 0.580 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.660 ;
END Via3_DV1N_eo

Via Via3_DV2E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.100 0.590 0.100 ;
    LAYER Via3 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.175 0.520 0.175 ;
END Via3_DV2E_eo

Via Via3_DV2EN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.100 0.590 0.180 ;
    LAYER Via3 ;
        RECT -0.090 -0.020 0.100 0.170 ;
        RECT  0.320 -0.020 0.510 0.170 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.250 ;
END Via3_DV2EN_eo

Via Via3_DV2ES_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.170 -0.180 0.590 0.100 ;
    LAYER Via3 ;
        RECT -0.090 -0.170 0.100 0.020 ;
        RECT  0.320 -0.170 0.510 0.020 ;
    LAYER Metal4 ;
        RECT -0.100 -0.250 0.520 0.100 ;
END Via3_DV2ES_eo

Via Via3_DV2W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.100  0.170 0.100 ;
    LAYER Via3 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal4 ;
        RECT -0.520 -0.175  0.100 0.175 ;
END Via3_DV2W_eo

Via Via3_DV2WN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.100  0.170 0.180 ;
    LAYER Via3 ;
        RECT -0.510 -0.020 -0.320 0.170 ;
        RECT -0.100 -0.020  0.090 0.170 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.250 ;
END Via3_DV2WN_eo

Via Via3_DV2WS_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.590 -0.180  0.170 0.100 ;
    LAYER Via3 ;
        RECT -0.510 -0.170 -0.320 0.020 ;
        RECT -0.100 -0.170  0.090 0.020 ;
    LAYER Metal4 ;
        RECT -0.520 -0.250  0.100 0.100 ;
END Via3_DV2WS_eo

Via Via3_DV2S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.175 -0.520 0.175  0.100 ;
    LAYER Via3 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.590 0.100  0.170 ;
END Via3_DV2S_eo

Via Via3_DV2SE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.520 0.250  0.100 ;
    LAYER Via3 ;
        RECT -0.020 -0.100 0.170  0.090 ;
        RECT -0.020 -0.510 0.170 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.590 0.220  0.170 ;
END Via3_DV2SE_eo

Via Via3_DV2SW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.520 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.170 -0.100 0.020  0.090 ;
        RECT -0.170 -0.510 0.020 -0.320 ;
    LAYER Metal4 ;
        RECT -0.220 -0.590 0.100  0.170 ;
END Via3_DV2SW_eo

Via Via3_DV2N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.175 -0.100 0.175 0.520 ;
    LAYER Via3 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.170 0.100 0.590 ;
END Via3_DV2N_eo

Via Via3_DV2NE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.250 0.520 ;
    LAYER Via3 ;
        RECT -0.020 -0.090 0.170 0.100 ;
        RECT -0.020  0.320 0.170 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.170 0.220 0.590 ;
END Via3_DV2NE_eo

Via Via3_DV2NW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.250 -0.100 0.100 0.520 ;
    LAYER Via3 ;
        RECT -0.170 -0.090 0.020 0.100 ;
        RECT -0.170  0.320 0.020 0.510 ;
    LAYER Metal4 ;
        RECT -0.220 -0.170 0.100 0.590 ;
END Via3_DV2NW_eo

##############

Via Via3_DV1EN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.100 0.660 0.190 ;
    LAYER Via3 ;
        RECT -0.020 -0.050 0.170 0.140 ;
        RECT  0.390 -0.050 0.580 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.660 0.190 ;
END Via3_DV1EN_beo

Via Via3_DV1ES_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.190 0.660 0.100 ;
    LAYER Via3 ;
        RECT -0.020 -0.140 0.170 0.050 ;
        RECT  0.390 -0.140 0.580 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.660 0.100 ;
END Via3_DV1ES_beo

Via Via3_DV1WN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.100  0.100 0.190 ;
    LAYER Via3 ;
        RECT -0.580 -0.050 -0.390 0.140 ;
        RECT -0.170 -0.050  0.020 0.140 ;
    LAYER Metal4 ;
        RECT -0.660 -0.100  0.100 0.190 ;
END Via3_DV1WN_beo

Via Via3_DV1WS_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.660 -0.190  0.100 0.100 ;
    LAYER Via3 ;
        RECT -0.580 -0.140 -0.390 0.050 ;
        RECT -0.170 -0.140  0.020 0.050 ;
    LAYER Metal4 ;
        RECT -0.660 -0.190  0.100 0.100 ;
END Via3_DV1WS_beo

Via Via3_DV1SE_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.100 -0.660 0.190  0.100 ;
    LAYER Via3 ;
        RECT -0.050 -0.170 0.140  0.020 ;
        RECT -0.050 -0.580 0.140 -0.390 ;
    LAYER Metal4 ;
        RECT -0.100 -0.660 0.190  0.100 ;
END Via3_DV1SE_beo

Via Via3_DV1SW_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal3 ;
        RECT -0.190 -0.660 0.100  0.100 ;
    LAYER Via3 ;
        RECT -0.140 -0.170 0.050  0.020 ;
        RECT -0.140 -0.580 0.050 -0.390 ;
    LAYER Metal4 ;
        RECT -0.190 -0.660 0.100  0.100 ;
END Via3_DV1SW_beo

Via Via4_XX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via4_XX_so

Via Via4_XXE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.190 0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.095 0.140 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.100 ;
END Via4_XXE_so

Via Via4_XXW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.100 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.095 0.050 0.095 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.100 ;
END Via4_XXW_so

Via Via4_YY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via4 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via4_YY_so

Via Via4_YYN_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.100 0.190 ;
    LAYER Via4 ;
        RECT -0.095 -0.050 0.095 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.190 ;
END Via4_YYN_so

Via Via4_YYS_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.190 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.140 0.095 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.100 0.100 ;
END Via4_YYS_so

Via Via4_XY_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.100 0.145 0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.100 0.145 ;
END Via4_XY_so

Via Via4_XYNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.100 0.100 0.150 ;
    LAYER Via4 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.150 -0.100 0.100 0.190 ;
END Via4_XYNW_so

Via Via4_XYNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.190 0.150 ;
    LAYER Via4 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.150 0.190 ;
END Via4_XYNE_so

Via Via4_XYSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.150 0.190 0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.150 0.100 ;
END Via4_XYSE_so

Via Via4_XYSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.150 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.150 -0.190 0.100 0.100 ;
END Via4_XYSW_so

Via Via4_YX_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.145 0.100 0.145 ;
    LAYER Via4 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.100 ;
END Via4_YX_so

Via Via4_YXNW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.150 -0.100 0.100 0.190 ;
    LAYER Via4 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.150 ;
END Via4_YXNW_so

Via Via4_YXNE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.150 0.190 ;
    LAYER Via4 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.150 ;
END Via4_YXNE_so

Via Via4_YXSE_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.190 0.150 0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.150 0.190 0.100 ;
END Via4_YXSE_so

Via Via4_YXSW_so DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.150 -0.190 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.190 -0.150 0.100 0.100 ;
END Via4_YXSW_so

##############

Via Via4_NE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.190 0.190 ;
    LAYER Via4 ;
        RECT -0.050 -0.050 0.140 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.190 ;
END Via4_NE_eo

Via Via4_NW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.100 0.100 0.190 ;
    LAYER Via4 ;
        RECT -0.140 -0.050 0.050 0.140 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.190 ;
END Via4_NW_eo

Via Via4_SE_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.190 0.190 0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.140 0.140 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.190 0.100 ;
END Via4_SE_eo

Via Via4_SW_eo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.190 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.140 0.050 0.050 ;
    LAYER Metal4 ;
        RECT -0.190 -0.190 0.100 0.100 ;
END Via4_SW_eo

##############

Via Via4_NE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.250 0.250 ;
    LAYER Via4 ;
        RECT -0.020 -0.020 0.170 0.170 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.250 0.250 ;
END Via4_NE_beo

Via Via4_NW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.250 -0.100 0.100 0.250 ;
    LAYER Via4 ;
        RECT -0.170 -0.020 0.020 0.170 ;
    LAYER Metal4 ;
        RECT -0.250 -0.100 0.100 0.250 ;
END Via4_NW_beo

Via Via4_SE_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.250 0.250 0.100 ;
    LAYER Via4 ;
        RECT -0.020 -0.170 0.170 0.020 ;
    LAYER Metal4 ;
        RECT -0.100 -0.250 0.250 0.100 ;
END Via4_SE_beo

Via Via4_SW_beo DEFAULT
    RESISTANCE 20.0 ;
    LAYER Metal5 ;
        RECT -0.250 -0.250 0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.170 -0.170 0.020 0.020 ;
    LAYER Metal4 ;
        RECT -0.250 -0.250 0.100 0.100 ;
END Via4_SW_beo

##############

Via Via4_DV1E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.600 0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.095 0.140 0.095 ;
        RECT  0.360 -0.095 0.550 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.600 0.100 ;
END Via4_DV1E_so

Via Via4_DV1W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.600 -0.100  0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.550 -0.095 -0.360 0.095 ;
        RECT -0.140 -0.095  0.050 0.095 ;
    LAYER Metal4 ;
        RECT -0.600 -0.100  0.100 0.100 ;
END Via4_DV1W_so

Via Via4_DV1S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.600 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.140 0.095  0.050 ;
        RECT -0.095 -0.550 0.095 -0.360 ;
    LAYER Metal4 ;
        RECT -0.100 -0.600 0.100  0.100 ;
END Via4_DV1S_so

Via Via4_DV1N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.100 0.600 ;
    LAYER Via4 ;
        RECT -0.095 -0.050 0.095 0.140 ;
        RECT -0.095  0.360 0.095 0.550 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.600 ;
END Via4_DV1N_so

Via Via4_DV2E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.140 -0.100 0.560 0.100 ;
    LAYER Via4 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via4_DV2E_so

Via Via4_DV2EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.140 -0.100 0.560 0.150 ;
    LAYER Via4 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via4_DV2EN_so

Via Via4_DV2ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.140 -0.150 0.560 0.100 ;
    LAYER Via4 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via4_DV2ES_so

Via Via4_DV2W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.560 -0.100  0.140 0.100 ;
    LAYER Via4 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal4 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via4_DV2W_so

Via Via4_DV2WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.560 -0.100  0.140 0.150 ;
    LAYER Via4 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via4_DV2WN_so

Via Via4_DV2WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.560 -0.150  0.140 0.100 ;
    LAYER Via4 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal4 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via4_DV2WS_so

Via Via4_DV2S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.560 0.100  0.140 ;
END Via4_DV2S_so

Via Via4_DV2SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.560 0.150  0.140 ;
END Via4_DV2SE_so

Via Via4_DV2SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal4 ;
        RECT -0.150 -0.560 0.100  0.140 ;
END Via4_DV2SW_so

Via Via4_DV2N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via4 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.140 0.100 0.560 ;
END Via4_DV2N_so

Via Via4_DV2NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via4 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.140 0.150 0.560 ;
END Via4_DV2NE_so

Via Via4_DV2NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via4 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal4 ;
        RECT -0.150 -0.140 0.100 0.560 ;
END Via4_DV2NW_so

##############

Via Via4_DV3E_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.145 0.520 0.145 ;
    LAYER Via4 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.145 0.520 0.145 ;
END Via4_DV3E_so

Via Via4_DV3EN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.520 0.190 ;
    LAYER Via4 ;
        RECT -0.090 -0.050 0.100 0.140 ;
        RECT  0.320 -0.050 0.510 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.190 ;
END Via4_DV3EN_so

Via Via4_DV3ES_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.190 0.520 0.100 ;
    LAYER Via4 ;
        RECT -0.090 -0.140 0.100 0.050 ;
        RECT  0.320 -0.140 0.510 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.520 0.100 ;
END Via4_DV3ES_so

Via Via4_DV3W_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.520 -0.145  0.100 0.145 ;
    LAYER Via4 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal4 ;
        RECT -0.520 -0.145  0.100 0.145 ;
END Via4_DV3W_so

Via Via4_DV3WN_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.520 -0.100  0.100 0.190 ;
    LAYER Via4 ;
        RECT -0.510 -0.050 -0.320 0.140 ;
        RECT -0.100 -0.050  0.090 0.140 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.190 ;
END Via4_DV3WN_so

Via Via4_DV3WS_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.520 -0.190  0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.510 -0.140 -0.320 0.050 ;
        RECT -0.100 -0.140  0.090 0.050 ;
    LAYER Metal4 ;
        RECT -0.520 -0.190  0.100 0.100 ;
END Via4_DV3WS_so

Via Via4_DV3S_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.520 0.145  0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal4 ;
        RECT -0.145 -0.520 0.145  0.100 ;
END Via4_DV3S_so

Via Via4_DV3SE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.520 0.190  0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.100 0.140  0.090 ;
        RECT -0.050 -0.510 0.140 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.520 0.190  0.100 ;
END Via4_DV3SE_so

Via Via4_DV3SW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.520 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.100 0.050  0.090 ;
        RECT -0.140 -0.510 0.050 -0.320 ;
    LAYER Metal4 ;
        RECT -0.190 -0.520 0.100  0.100 ;
END Via4_DV3SW_so

Via Via4_DV3N_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.145 -0.100 0.145 0.520 ;
    LAYER Via4 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal4 ;
        RECT -0.145 -0.100 0.145 0.520 ;
END Via4_DV3N_so

Via Via4_DV3NE_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.190 0.520 ;
    LAYER Via4 ;
        RECT -0.050 -0.090 0.140 0.100 ;
        RECT -0.050  0.320 0.140 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.190 0.520 ;
END Via4_DV3NE_so

Via Via4_DV3NW_so DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.100 0.100 0.520 ;
    LAYER Via4 ;
        RECT -0.140 -0.090 0.050 0.100 ;
        RECT -0.140  0.320 0.050 0.510 ;
    LAYER Metal4 ;
        RECT -0.190 -0.100 0.100 0.520 ;
END Via4_DV3NW_so

##############

Via Via4_DV1E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.660 0.100 ;
    LAYER Via4 ;
        RECT -0.020 -0.095 0.170 0.095 ;
        RECT  0.390 -0.095 0.580 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.660 0.100 ;
END Via4_DV1E_eo

Via Via4_DV1W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.660 -0.100  0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.580 -0.095 -0.390 0.095 ;
        RECT -0.170 -0.095  0.020 0.095 ;
    LAYER Metal4 ;
        RECT -0.660 -0.100  0.100 0.100 ;
END Via4_DV1W_eo

Via Via4_DV1S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.660 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.170 0.095  0.020 ;
        RECT -0.095 -0.580 0.095 -0.390 ;
    LAYER Metal4 ;
        RECT -0.100 -0.660 0.100  0.100 ;
END Via4_DV1S_eo

Via Via4_DV1N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.100 0.660 ;
    LAYER Via4 ;
        RECT -0.095 -0.020 0.095 0.170 ;
        RECT -0.095  0.390 0.095 0.580 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.100 0.660 ;
END Via4_DV1N_eo

Via Via4_DV2E_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.170 -0.100 0.590 0.100 ;
    LAYER Via4 ;
        RECT -0.090 -0.095 0.100 0.095 ;
        RECT  0.320 -0.095 0.510 0.095 ;
    LAYER Metal4 ;
        RECT -0.100 -0.175 0.520 0.175 ;
END Via4_DV2E_eo

Via Via4_DV2EN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.170 -0.100 0.590 0.180 ;
    LAYER Via4 ;
        RECT -0.090 -0.020 0.100 0.170 ;
        RECT  0.320 -0.020 0.510 0.170 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.520 0.250 ;
END Via4_DV2EN_eo

Via Via4_DV2ES_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.170 -0.180 0.590 0.100 ;
    LAYER Via4 ;
        RECT -0.090 -0.170 0.100 0.020 ;
        RECT  0.320 -0.170 0.510 0.020 ;
    LAYER Metal4 ;
        RECT -0.100 -0.250 0.520 0.100 ;
END Via4_DV2ES_eo

Via Via4_DV2W_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.590 -0.100  0.170 0.100 ;
    LAYER Via4 ;
        RECT -0.510 -0.095 -0.320 0.095 ;
        RECT -0.100 -0.095  0.090 0.095 ;
    LAYER Metal4 ;
        RECT -0.520 -0.175  0.100 0.175 ;
END Via4_DV2W_eo

Via Via4_DV2WN_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.590 -0.100  0.170 0.180 ;
    LAYER Via4 ;
        RECT -0.510 -0.020 -0.320 0.170 ;
        RECT -0.100 -0.020  0.090 0.170 ;
    LAYER Metal4 ;
        RECT -0.520 -0.100  0.100 0.250 ;
END Via4_DV2WN_eo

Via Via4_DV2WS_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.590 -0.180  0.170 0.100 ;
    LAYER Via4 ;
        RECT -0.510 -0.170 -0.320 0.020 ;
        RECT -0.100 -0.170  0.090 0.020 ;
    LAYER Metal4 ;
        RECT -0.520 -0.250  0.100 0.100 ;
END Via4_DV2WS_eo

Via Via4_DV2S_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.175 -0.520 0.175  0.100 ;
    LAYER Via4 ;
        RECT -0.095 -0.100 0.095  0.090 ;
        RECT -0.095 -0.510 0.095 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.590 0.100  0.170 ;
END Via4_DV2S_eo

Via Via4_DV2SE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.520 0.250  0.100 ;
    LAYER Via4 ;
        RECT -0.020 -0.100 0.170  0.090 ;
        RECT -0.020 -0.510 0.170 -0.320 ;
    LAYER Metal4 ;
        RECT -0.100 -0.590 0.220  0.170 ;
END Via4_DV2SE_eo

Via Via4_DV2SW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.250 -0.520 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.170 -0.100 0.020  0.090 ;
        RECT -0.170 -0.510 0.020 -0.320 ;
    LAYER Metal4 ;
        RECT -0.220 -0.590 0.100  0.170 ;
END Via4_DV2SW_eo

Via Via4_DV2N_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.175 -0.100 0.175 0.520 ;
    LAYER Via4 ;
        RECT -0.095 -0.090 0.095 0.100 ;
        RECT -0.095  0.320 0.095 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.170 0.100 0.590 ;
END Via4_DV2N_eo

Via Via4_DV2NE_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.250 0.520 ;
    LAYER Via4 ;
        RECT -0.020 -0.090 0.170 0.100 ;
        RECT -0.020  0.320 0.170 0.510 ;
    LAYER Metal4 ;
        RECT -0.100 -0.170 0.220 0.590 ;
END Via4_DV2NE_eo

Via Via4_DV2NW_eo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.250 -0.100 0.100 0.520 ;
    LAYER Via4 ;
        RECT -0.170 -0.090 0.020 0.100 ;
        RECT -0.170  0.320 0.020 0.510 ;
    LAYER Metal4 ;
        RECT -0.220 -0.170 0.100 0.590 ;
END Via4_DV2NW_eo

##############

Via Via4_DV1EN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.100 0.660 0.190 ;
    LAYER Via4 ;
        RECT -0.020 -0.050 0.170 0.140 ;
        RECT  0.390 -0.050 0.580 0.140 ;
    LAYER Metal4 ;
        RECT -0.100 -0.100 0.660 0.190 ;
END Via4_DV1EN_beo

Via Via4_DV1ES_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.190 0.660 0.100 ;
    LAYER Via4 ;
        RECT -0.020 -0.140 0.170 0.050 ;
        RECT  0.390 -0.140 0.580 0.050 ;
    LAYER Metal4 ;
        RECT -0.100 -0.190 0.660 0.100 ;
END Via4_DV1ES_beo

Via Via4_DV1WN_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.660 -0.100  0.100 0.190 ;
    LAYER Via4 ;
        RECT -0.580 -0.050 -0.390 0.140 ;
        RECT -0.170 -0.050  0.020 0.140 ;
    LAYER Metal4 ;
        RECT -0.660 -0.100  0.100 0.190 ;
END Via4_DV1WN_beo

Via Via4_DV1WS_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.660 -0.190  0.100 0.100 ;
    LAYER Via4 ;
        RECT -0.580 -0.140 -0.390 0.050 ;
        RECT -0.170 -0.140  0.020 0.050 ;
    LAYER Metal4 ;
        RECT -0.660 -0.190  0.100 0.100 ;
END Via4_DV1WS_beo

Via Via4_DV1SE_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.100 -0.660 0.190  0.100 ;
    LAYER Via4 ;
        RECT -0.050 -0.170 0.140  0.020 ;
        RECT -0.050 -0.580 0.140 -0.390 ;
    LAYER Metal4 ;
        RECT -0.100 -0.660 0.190  0.100 ;
END Via4_DV1SE_beo

Via Via4_DV1SW_beo DEFAULT
    RESISTANCE 10.0 ;
    LAYER Metal5 ;
        RECT -0.190 -0.660 0.100  0.100 ;
    LAYER Via4 ;
        RECT -0.140 -0.170 0.050  0.020 ;
        RECT -0.140 -0.580 0.050 -0.390 ;
    LAYER Metal4 ;
        RECT -0.190 -0.660 0.100  0.100 ;
END Via4_DV1SW_beo
########################################
Via TopVia1EWNS DEFAULT
  RESISTANCE 4.0 ;
  LAYER Metal5 ;
    RECT -0.31 -0.31 0.31 0.31 ;
  LAYER TopVia1 ;
    RECT -0.21 -0.21 0.21 0.21 ;
  LAYER TopMetal1 ;
    RECT -0.75 -0.75 0.75 0.75 ;
END TopVia1EWNS

Via TopVia2EWNS DEFAULT
  RESISTANCE 2.2 ;
  LAYER TopMetal1 ;
    RECT -0.95 -0.95 0.95 0.95 ;
  LAYER TopVia2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
  LAYER TopMetal2 ;
    RECT -0.95 -0.95 0.95 0.95 ;
END TopVia2EWNS
#########################################
ViaRULE via1Array GENERATE
    LAYER Metal1 ;
        ENCLOSURE 0.050 0.010 ;

    LAYER Metal2 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Via1 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
        RESISTANCE 20.0 ;
END via1Array

ViaRULE via2Array GENERATE
    LAYER Metal2 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Metal3 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Via2 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
        RESISTANCE 20.0 ;
END via2Array

ViaRULE via3Array GENERATE
    LAYER Metal3 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Metal4 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Via3 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
        RESISTANCE 20.0 ;
END via3Array

ViaRULE via4Array GENERATE
    LAYER Metal4 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Metal5 ;
        ENCLOSURE 0.050 0.005 ;

    LAYER Via4 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
        RESISTANCE 20.0 ;
END via4Array
###########################################
ViaRULE viagen56 GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0 0 ;
  LAYER TopMetal1 ;
    ENCLOSURE 0.61 0.61 ;
  LAYER TopVia1 ;
    RECT -0.21 -0.21 0.21 0.21 ;
    SPACING 0.84 BY 0.84 ;
    RESISTANCE 4.0 ;
END viagen56

ViaRULE viagen67 GENERATE
  LAYER TopMetal1 ;
    ENCLOSURE 0.5 0.5 ;
  LAYER TopMetal2 ;
    ENCLOSURE 0.55 0.55 ;
  LAYER TopVia2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
    SPACING 1.96 BY 1.96 ;
    RESISTANCE 2.2 ;
END viagen67

END LIBRARY

